/* External Modules
module test_pe (
  input  bit0,
  input  bit1,
  input  bit2,
  input [7:0] cfg_a,
  input [31:0] cfg_d,
  input  cfg_en,
  input  clk,
  input  clk_en,
  input [15:0] data0,
  input [15:0] data1,
  output  irq,
  output [31:0] read_data,
  output [15:0] res,
  output  res_p,
  input  rst_n
);

endmodule  // test_pe

*/
module coreir_ult #(parameter width=1) (
  input [width-1:0] in0,
  input [width-1:0] in1,
  output out
);
  assign out = in0 < in1;

endmodule  // coreir_ult

module coreir_slice #(parameter hi=1, parameter lo=0, parameter width=1) (
  input [width-1:0] in,
  output [hi-lo-1:0] out
);
  assign out = in[hi-1:lo];

endmodule  // coreir_slice

module coreir_reg_arst #(parameter arst_posedge=1, parameter clk_posedge=1, parameter init=1, parameter width=1) (
  input clk,
  input arst,
  input [width-1:0] in,
  output [width-1:0] out
);
  reg [width-1:0] outReg;
  wire real_rst;
  assign real_rst = arst_posedge ? arst : ~arst;
  wire real_clk;
  assign real_clk = clk_posedge ? clk : ~clk;
  always @(posedge real_clk, posedge real_rst) begin
    if (real_rst) outReg <= init;
    else outReg <= in;
  end
  assign out = outReg;

endmodule  // coreir_reg_arst

module coreir_reg #(parameter clk_posedge=1, parameter init=1, parameter width=1) (
  input clk,
  input [width-1:0] in,
  output [width-1:0] out
);
  reg [width-1:0] outReg=init;
  wire real_clk;
  assign real_clk = clk_posedge ? clk : ~clk;
  always @(posedge real_clk) begin
    outReg <= in;
  end
  assign out = outReg;

endmodule  // coreir_reg

module coreir_not #(parameter width=1) (
  input [width-1:0] in,
  output [width-1:0] out
);
  assign out = ~in;

endmodule  // coreir_not

module coreir_mux #(parameter width=1) (
  input [width-1:0] in0,
  input [width-1:0] in1,
  input sel,
  output [width-1:0] out
);
  assign out = sel ? in1 : in0;

endmodule  // coreir_mux

module coreir_eq #(parameter width=1) (
  input [width-1:0] in0,
  input [width-1:0] in1,
  output out
);
  assign out = in0 == in1;

endmodule  // coreir_eq

module coreir_const #(parameter value=1, parameter width=1) (
  output [width-1:0] out
);
  assign out = value;

endmodule  // coreir_const

module corebit_term (
  input in
);


endmodule  // corebit_term

module corebit_const #(parameter value=1) (
  output out
);
  assign out = value;

endmodule  // corebit_const

module corebit_and (
  input in0,
  input in1,
  output out
);
  assign out = in0 & in1;

endmodule  // corebit_and

// Generated from commonlib.muxn(N:2, width:4)
module commonlib_muxn__N2__width4 (
  input [3:0] in_data_0,
  input [3:0] in_data_1,
  input [0:0] in_sel,
  output [3:0] out
);


  // Instancing generated Module: coreir.mux(width:4)
  wire [3:0] _join__in0;
  wire [3:0] _join__in1;
  wire [3:0] _join__out;
  wire  _join__sel;
  coreir_mux #(.width(4)) _join(
    .in0(_join__in0),
    .in1(_join__in1),
    .out(_join__out),
    .sel(_join__sel)
  );

  assign _join__in0[3:0] = in_data_0[3:0];

  assign _join__in1[3:0] = in_data_1[3:0];

  assign out[3:0] = _join__out[3:0];

  assign _join__sel = in_sel[0];


endmodule  // commonlib_muxn__N2__width4

// Generated from commonlib.muxn(N:2, width:32)
module commonlib_muxn__N2__width32 (
  input [31:0] in_data_0,
  input [31:0] in_data_1,
  input [0:0] in_sel,
  output [31:0] out
);


  // Instancing generated Module: coreir.mux(width:32)
  wire [31:0] _join__in0;
  wire [31:0] _join__in1;
  wire [31:0] _join__out;
  wire  _join__sel;
  coreir_mux #(.width(32)) _join(
    .in0(_join__in0),
    .in1(_join__in1),
    .out(_join__out),
    .sel(_join__sel)
  );

  assign _join__in0[31:0] = in_data_0[31:0];

  assign _join__in1[31:0] = in_data_1[31:0];

  assign out[31:0] = _join__out[31:0];

  assign _join__sel = in_sel[0];


endmodule  // commonlib_muxn__N2__width32

// Generated from commonlib.muxn(N:4, width:32)
module commonlib_muxn__N4__width32 (
  input [31:0] in_data_0,
  input [31:0] in_data_1,
  input [31:0] in_data_2,
  input [31:0] in_data_3,
  input [1:0] in_sel,
  output [31:0] out
);


  // Instancing generated Module: coreir.mux(width:32)
  wire [31:0] _join__in0;
  wire [31:0] _join__in1;
  wire [31:0] _join__out;
  wire  _join__sel;
  coreir_mux #(.width(32)) _join(
    .in0(_join__in0),
    .in1(_join__in1),
    .out(_join__out),
    .sel(_join__sel)
  );

  // Instancing generated Module: commonlib.muxn(N:2, width:32)
  wire [31:0] muxN_0__in_data_0;
  wire [31:0] muxN_0__in_data_1;
  wire [0:0] muxN_0__in_sel;
  wire [31:0] muxN_0__out;
  commonlib_muxn__N2__width32 muxN_0(
    .in_data_0(muxN_0__in_data_0),
    .in_data_1(muxN_0__in_data_1),
    .in_sel(muxN_0__in_sel),
    .out(muxN_0__out)
  );

  // Instancing generated Module: commonlib.muxn(N:2, width:32)
  wire [31:0] muxN_1__in_data_0;
  wire [31:0] muxN_1__in_data_1;
  wire [0:0] muxN_1__in_sel;
  wire [31:0] muxN_1__out;
  commonlib_muxn__N2__width32 muxN_1(
    .in_data_0(muxN_1__in_data_0),
    .in_data_1(muxN_1__in_data_1),
    .in_sel(muxN_1__in_sel),
    .out(muxN_1__out)
  );

  // Instancing generated Module: coreir.slice(hi:1, lo:0, width:2)
  wire [1:0] sel_slice0__in;
  wire [0:0] sel_slice0__out;
  coreir_slice #(.hi(1),.lo(0),.width(2)) sel_slice0(
    .in(sel_slice0__in),
    .out(sel_slice0__out)
  );

  // Instancing generated Module: coreir.slice(hi:1, lo:0, width:2)
  wire [1:0] sel_slice1__in;
  wire [0:0] sel_slice1__out;
  coreir_slice #(.hi(1),.lo(0),.width(2)) sel_slice1(
    .in(sel_slice1__in),
    .out(sel_slice1__out)
  );

  assign _join__in0[31:0] = muxN_0__out[31:0];

  assign _join__in1[31:0] = muxN_1__out[31:0];

  assign out[31:0] = _join__out[31:0];

  assign _join__sel = in_sel[1];

  assign muxN_0__in_data_0[31:0] = in_data_0[31:0];

  assign muxN_0__in_data_1[31:0] = in_data_1[31:0];

  assign muxN_0__in_sel[0:0] = sel_slice0__out[0:0];

  assign muxN_1__in_data_0[31:0] = in_data_2[31:0];

  assign muxN_1__in_data_1[31:0] = in_data_3[31:0];

  assign muxN_1__in_sel[0:0] = sel_slice1__out[0:0];

  assign sel_slice0__in[1:0] = in_sel[1:0];

  assign sel_slice1__in[1:0] = in_sel[1:0];


endmodule  // commonlib_muxn__N4__width32

// Generated from commonlib.muxn(N:8, width:32)
module commonlib_muxn__N8__width32 (
  input [31:0] in_data_0,
  input [31:0] in_data_1,
  input [31:0] in_data_2,
  input [31:0] in_data_3,
  input [31:0] in_data_4,
  input [31:0] in_data_5,
  input [31:0] in_data_6,
  input [31:0] in_data_7,
  input [2:0] in_sel,
  output [31:0] out
);


  // Instancing generated Module: coreir.mux(width:32)
  wire [31:0] _join__in0;
  wire [31:0] _join__in1;
  wire [31:0] _join__out;
  wire  _join__sel;
  coreir_mux #(.width(32)) _join(
    .in0(_join__in0),
    .in1(_join__in1),
    .out(_join__out),
    .sel(_join__sel)
  );

  // Instancing generated Module: commonlib.muxn(N:4, width:32)
  wire [31:0] muxN_0__in_data_0;
  wire [31:0] muxN_0__in_data_1;
  wire [31:0] muxN_0__in_data_2;
  wire [31:0] muxN_0__in_data_3;
  wire [1:0] muxN_0__in_sel;
  wire [31:0] muxN_0__out;
  commonlib_muxn__N4__width32 muxN_0(
    .in_data_0(muxN_0__in_data_0),
    .in_data_1(muxN_0__in_data_1),
    .in_data_2(muxN_0__in_data_2),
    .in_data_3(muxN_0__in_data_3),
    .in_sel(muxN_0__in_sel),
    .out(muxN_0__out)
  );

  // Instancing generated Module: commonlib.muxn(N:4, width:32)
  wire [31:0] muxN_1__in_data_0;
  wire [31:0] muxN_1__in_data_1;
  wire [31:0] muxN_1__in_data_2;
  wire [31:0] muxN_1__in_data_3;
  wire [1:0] muxN_1__in_sel;
  wire [31:0] muxN_1__out;
  commonlib_muxn__N4__width32 muxN_1(
    .in_data_0(muxN_1__in_data_0),
    .in_data_1(muxN_1__in_data_1),
    .in_data_2(muxN_1__in_data_2),
    .in_data_3(muxN_1__in_data_3),
    .in_sel(muxN_1__in_sel),
    .out(muxN_1__out)
  );

  // Instancing generated Module: coreir.slice(hi:2, lo:0, width:3)
  wire [2:0] sel_slice0__in;
  wire [1:0] sel_slice0__out;
  coreir_slice #(.hi(2),.lo(0),.width(3)) sel_slice0(
    .in(sel_slice0__in),
    .out(sel_slice0__out)
  );

  // Instancing generated Module: coreir.slice(hi:2, lo:0, width:3)
  wire [2:0] sel_slice1__in;
  wire [1:0] sel_slice1__out;
  coreir_slice #(.hi(2),.lo(0),.width(3)) sel_slice1(
    .in(sel_slice1__in),
    .out(sel_slice1__out)
  );

  assign _join__in0[31:0] = muxN_0__out[31:0];

  assign _join__in1[31:0] = muxN_1__out[31:0];

  assign out[31:0] = _join__out[31:0];

  assign _join__sel = in_sel[2];

  assign muxN_0__in_data_0[31:0] = in_data_0[31:0];

  assign muxN_0__in_data_1[31:0] = in_data_1[31:0];

  assign muxN_0__in_data_2[31:0] = in_data_2[31:0];

  assign muxN_0__in_data_3[31:0] = in_data_3[31:0];

  assign muxN_0__in_sel[1:0] = sel_slice0__out[1:0];

  assign muxN_1__in_data_0[31:0] = in_data_4[31:0];

  assign muxN_1__in_data_1[31:0] = in_data_5[31:0];

  assign muxN_1__in_data_2[31:0] = in_data_6[31:0];

  assign muxN_1__in_data_3[31:0] = in_data_7[31:0];

  assign muxN_1__in_sel[1:0] = sel_slice1__out[1:0];

  assign sel_slice0__in[2:0] = in_sel[2:0];

  assign sel_slice1__in[2:0] = in_sel[2:0];


endmodule  // commonlib_muxn__N8__width32

// Generated from commonlib.muxn(N:2, width:2)
module commonlib_muxn__N2__width2 (
  input [1:0] in_data_0,
  input [1:0] in_data_1,
  input [0:0] in_sel,
  output [1:0] out
);


  // Instancing generated Module: coreir.mux(width:2)
  wire [1:0] _join__in0;
  wire [1:0] _join__in1;
  wire [1:0] _join__out;
  wire  _join__sel;
  coreir_mux #(.width(2)) _join(
    .in0(_join__in0),
    .in1(_join__in1),
    .out(_join__out),
    .sel(_join__sel)
  );

  assign _join__in0[1:0] = in_data_0[1:0];

  assign _join__in1[1:0] = in_data_1[1:0];

  assign out[1:0] = _join__out[1:0];

  assign _join__sel = in_sel[0];


endmodule  // commonlib_muxn__N2__width2

// Generated from commonlib.muxn(N:2, width:16)
module commonlib_muxn__N2__width16 (
  input [15:0] in_data_0,
  input [15:0] in_data_1,
  input [0:0] in_sel,
  output [15:0] out
);


  // Instancing generated Module: coreir.mux(width:16)
  wire [15:0] _join__in0;
  wire [15:0] _join__in1;
  wire [15:0] _join__out;
  wire  _join__sel;
  coreir_mux #(.width(16)) _join(
    .in0(_join__in0),
    .in1(_join__in1),
    .out(_join__out),
    .sel(_join__sel)
  );

  assign _join__in0[15:0] = in_data_0[15:0];

  assign _join__in1[15:0] = in_data_1[15:0];

  assign out[15:0] = _join__out[15:0];

  assign _join__sel = in_sel[0];


endmodule  // commonlib_muxn__N2__width16

// Generated from commonlib.muxn(N:4, width:16)
module commonlib_muxn__N4__width16 (
  input [15:0] in_data_0,
  input [15:0] in_data_1,
  input [15:0] in_data_2,
  input [15:0] in_data_3,
  input [1:0] in_sel,
  output [15:0] out
);


  // Instancing generated Module: coreir.mux(width:16)
  wire [15:0] _join__in0;
  wire [15:0] _join__in1;
  wire [15:0] _join__out;
  wire  _join__sel;
  coreir_mux #(.width(16)) _join(
    .in0(_join__in0),
    .in1(_join__in1),
    .out(_join__out),
    .sel(_join__sel)
  );

  // Instancing generated Module: commonlib.muxn(N:2, width:16)
  wire [15:0] muxN_0__in_data_0;
  wire [15:0] muxN_0__in_data_1;
  wire [0:0] muxN_0__in_sel;
  wire [15:0] muxN_0__out;
  commonlib_muxn__N2__width16 muxN_0(
    .in_data_0(muxN_0__in_data_0),
    .in_data_1(muxN_0__in_data_1),
    .in_sel(muxN_0__in_sel),
    .out(muxN_0__out)
  );

  // Instancing generated Module: commonlib.muxn(N:2, width:16)
  wire [15:0] muxN_1__in_data_0;
  wire [15:0] muxN_1__in_data_1;
  wire [0:0] muxN_1__in_sel;
  wire [15:0] muxN_1__out;
  commonlib_muxn__N2__width16 muxN_1(
    .in_data_0(muxN_1__in_data_0),
    .in_data_1(muxN_1__in_data_1),
    .in_sel(muxN_1__in_sel),
    .out(muxN_1__out)
  );

  // Instancing generated Module: coreir.slice(hi:1, lo:0, width:2)
  wire [1:0] sel_slice0__in;
  wire [0:0] sel_slice0__out;
  coreir_slice #(.hi(1),.lo(0),.width(2)) sel_slice0(
    .in(sel_slice0__in),
    .out(sel_slice0__out)
  );

  // Instancing generated Module: coreir.slice(hi:1, lo:0, width:2)
  wire [1:0] sel_slice1__in;
  wire [0:0] sel_slice1__out;
  coreir_slice #(.hi(1),.lo(0),.width(2)) sel_slice1(
    .in(sel_slice1__in),
    .out(sel_slice1__out)
  );

  assign _join__in0[15:0] = muxN_0__out[15:0];

  assign _join__in1[15:0] = muxN_1__out[15:0];

  assign out[15:0] = _join__out[15:0];

  assign _join__sel = in_sel[1];

  assign muxN_0__in_data_0[15:0] = in_data_0[15:0];

  assign muxN_0__in_data_1[15:0] = in_data_1[15:0];

  assign muxN_0__in_sel[0:0] = sel_slice0__out[0:0];

  assign muxN_1__in_data_0[15:0] = in_data_2[15:0];

  assign muxN_1__in_data_1[15:0] = in_data_3[15:0];

  assign muxN_1__in_sel[0:0] = sel_slice1__out[0:0];

  assign sel_slice0__in[1:0] = in_sel[1:0];

  assign sel_slice1__in[1:0] = in_sel[1:0];


endmodule  // commonlib_muxn__N4__width16

// Generated from commonlib.muxn(N:8, width:16)
module commonlib_muxn__N8__width16 (
  input [15:0] in_data_0,
  input [15:0] in_data_1,
  input [15:0] in_data_2,
  input [15:0] in_data_3,
  input [15:0] in_data_4,
  input [15:0] in_data_5,
  input [15:0] in_data_6,
  input [15:0] in_data_7,
  input [2:0] in_sel,
  output [15:0] out
);


  // Instancing generated Module: coreir.mux(width:16)
  wire [15:0] _join__in0;
  wire [15:0] _join__in1;
  wire [15:0] _join__out;
  wire  _join__sel;
  coreir_mux #(.width(16)) _join(
    .in0(_join__in0),
    .in1(_join__in1),
    .out(_join__out),
    .sel(_join__sel)
  );

  // Instancing generated Module: commonlib.muxn(N:4, width:16)
  wire [15:0] muxN_0__in_data_0;
  wire [15:0] muxN_0__in_data_1;
  wire [15:0] muxN_0__in_data_2;
  wire [15:0] muxN_0__in_data_3;
  wire [1:0] muxN_0__in_sel;
  wire [15:0] muxN_0__out;
  commonlib_muxn__N4__width16 muxN_0(
    .in_data_0(muxN_0__in_data_0),
    .in_data_1(muxN_0__in_data_1),
    .in_data_2(muxN_0__in_data_2),
    .in_data_3(muxN_0__in_data_3),
    .in_sel(muxN_0__in_sel),
    .out(muxN_0__out)
  );

  // Instancing generated Module: commonlib.muxn(N:4, width:16)
  wire [15:0] muxN_1__in_data_0;
  wire [15:0] muxN_1__in_data_1;
  wire [15:0] muxN_1__in_data_2;
  wire [15:0] muxN_1__in_data_3;
  wire [1:0] muxN_1__in_sel;
  wire [15:0] muxN_1__out;
  commonlib_muxn__N4__width16 muxN_1(
    .in_data_0(muxN_1__in_data_0),
    .in_data_1(muxN_1__in_data_1),
    .in_data_2(muxN_1__in_data_2),
    .in_data_3(muxN_1__in_data_3),
    .in_sel(muxN_1__in_sel),
    .out(muxN_1__out)
  );

  // Instancing generated Module: coreir.slice(hi:2, lo:0, width:3)
  wire [2:0] sel_slice0__in;
  wire [1:0] sel_slice0__out;
  coreir_slice #(.hi(2),.lo(0),.width(3)) sel_slice0(
    .in(sel_slice0__in),
    .out(sel_slice0__out)
  );

  // Instancing generated Module: coreir.slice(hi:2, lo:0, width:3)
  wire [2:0] sel_slice1__in;
  wire [1:0] sel_slice1__out;
  coreir_slice #(.hi(2),.lo(0),.width(3)) sel_slice1(
    .in(sel_slice1__in),
    .out(sel_slice1__out)
  );

  assign _join__in0[15:0] = muxN_0__out[15:0];

  assign _join__in1[15:0] = muxN_1__out[15:0];

  assign out[15:0] = _join__out[15:0];

  assign _join__sel = in_sel[2];

  assign muxN_0__in_data_0[15:0] = in_data_0[15:0];

  assign muxN_0__in_data_1[15:0] = in_data_1[15:0];

  assign muxN_0__in_data_2[15:0] = in_data_2[15:0];

  assign muxN_0__in_data_3[15:0] = in_data_3[15:0];

  assign muxN_0__in_sel[1:0] = sel_slice0__out[1:0];

  assign muxN_1__in_data_0[15:0] = in_data_4[15:0];

  assign muxN_1__in_data_1[15:0] = in_data_5[15:0];

  assign muxN_1__in_data_2[15:0] = in_data_6[15:0];

  assign muxN_1__in_data_3[15:0] = in_data_7[15:0];

  assign muxN_1__in_sel[1:0] = sel_slice1__out[1:0];

  assign sel_slice0__in[2:0] = in_sel[2:0];

  assign sel_slice1__in[2:0] = in_sel[2:0];


endmodule  // commonlib_muxn__N8__width16

// Generated from commonlib.muxn(N:2, width:1)
module commonlib_muxn__N2__width1 (
  input [0:0] in_data_0,
  input [0:0] in_data_1,
  input [0:0] in_sel,
  output [0:0] out
);


  // Instancing generated Module: coreir.mux(width:1)
  wire [0:0] _join__in0;
  wire [0:0] _join__in1;
  wire [0:0] _join__out;
  wire  _join__sel;
  coreir_mux #(.width(1)) _join(
    .in0(_join__in0),
    .in1(_join__in1),
    .out(_join__out),
    .sel(_join__sel)
  );

  assign _join__in0[0:0] = in_data_0[0:0];

  assign _join__in1[0:0] = in_data_1[0:0];

  assign out[0:0] = _join__out[0:0];

  assign _join__sel = in_sel[0];


endmodule  // commonlib_muxn__N2__width1

// Generated from commonlib.muxn(N:4, width:1)
module commonlib_muxn__N4__width1 (
  input [0:0] in_data_0,
  input [0:0] in_data_1,
  input [0:0] in_data_2,
  input [0:0] in_data_3,
  input [1:0] in_sel,
  output [0:0] out
);


  // Instancing generated Module: coreir.mux(width:1)
  wire [0:0] _join__in0;
  wire [0:0] _join__in1;
  wire [0:0] _join__out;
  wire  _join__sel;
  coreir_mux #(.width(1)) _join(
    .in0(_join__in0),
    .in1(_join__in1),
    .out(_join__out),
    .sel(_join__sel)
  );

  // Instancing generated Module: commonlib.muxn(N:2, width:1)
  wire [0:0] muxN_0__in_data_0;
  wire [0:0] muxN_0__in_data_1;
  wire [0:0] muxN_0__in_sel;
  wire [0:0] muxN_0__out;
  commonlib_muxn__N2__width1 muxN_0(
    .in_data_0(muxN_0__in_data_0),
    .in_data_1(muxN_0__in_data_1),
    .in_sel(muxN_0__in_sel),
    .out(muxN_0__out)
  );

  // Instancing generated Module: commonlib.muxn(N:2, width:1)
  wire [0:0] muxN_1__in_data_0;
  wire [0:0] muxN_1__in_data_1;
  wire [0:0] muxN_1__in_sel;
  wire [0:0] muxN_1__out;
  commonlib_muxn__N2__width1 muxN_1(
    .in_data_0(muxN_1__in_data_0),
    .in_data_1(muxN_1__in_data_1),
    .in_sel(muxN_1__in_sel),
    .out(muxN_1__out)
  );

  // Instancing generated Module: coreir.slice(hi:1, lo:0, width:2)
  wire [1:0] sel_slice0__in;
  wire [0:0] sel_slice0__out;
  coreir_slice #(.hi(1),.lo(0),.width(2)) sel_slice0(
    .in(sel_slice0__in),
    .out(sel_slice0__out)
  );

  // Instancing generated Module: coreir.slice(hi:1, lo:0, width:2)
  wire [1:0] sel_slice1__in;
  wire [0:0] sel_slice1__out;
  coreir_slice #(.hi(1),.lo(0),.width(2)) sel_slice1(
    .in(sel_slice1__in),
    .out(sel_slice1__out)
  );

  assign _join__in0[0:0] = muxN_0__out[0:0];

  assign _join__in1[0:0] = muxN_1__out[0:0];

  assign out[0:0] = _join__out[0:0];

  assign _join__sel = in_sel[1];

  assign muxN_0__in_data_0[0:0] = in_data_0[0:0];

  assign muxN_0__in_data_1[0:0] = in_data_1[0:0];

  assign muxN_0__in_sel[0:0] = sel_slice0__out[0:0];

  assign muxN_1__in_data_0[0:0] = in_data_2[0:0];

  assign muxN_1__in_data_1[0:0] = in_data_3[0:0];

  assign muxN_1__in_sel[0:0] = sel_slice1__out[0:0];

  assign sel_slice0__in[1:0] = in_sel[1:0];

  assign sel_slice1__in[1:0] = in_sel[1:0];


endmodule  // commonlib_muxn__N4__width1

// Generated from commonlib.muxn(N:8, width:1)
module commonlib_muxn__N8__width1 (
  input [0:0] in_data_0,
  input [0:0] in_data_1,
  input [0:0] in_data_2,
  input [0:0] in_data_3,
  input [0:0] in_data_4,
  input [0:0] in_data_5,
  input [0:0] in_data_6,
  input [0:0] in_data_7,
  input [2:0] in_sel,
  output [0:0] out
);


  // Instancing generated Module: coreir.mux(width:1)
  wire [0:0] _join__in0;
  wire [0:0] _join__in1;
  wire [0:0] _join__out;
  wire  _join__sel;
  coreir_mux #(.width(1)) _join(
    .in0(_join__in0),
    .in1(_join__in1),
    .out(_join__out),
    .sel(_join__sel)
  );

  // Instancing generated Module: commonlib.muxn(N:4, width:1)
  wire [0:0] muxN_0__in_data_0;
  wire [0:0] muxN_0__in_data_1;
  wire [0:0] muxN_0__in_data_2;
  wire [0:0] muxN_0__in_data_3;
  wire [1:0] muxN_0__in_sel;
  wire [0:0] muxN_0__out;
  commonlib_muxn__N4__width1 muxN_0(
    .in_data_0(muxN_0__in_data_0),
    .in_data_1(muxN_0__in_data_1),
    .in_data_2(muxN_0__in_data_2),
    .in_data_3(muxN_0__in_data_3),
    .in_sel(muxN_0__in_sel),
    .out(muxN_0__out)
  );

  // Instancing generated Module: commonlib.muxn(N:4, width:1)
  wire [0:0] muxN_1__in_data_0;
  wire [0:0] muxN_1__in_data_1;
  wire [0:0] muxN_1__in_data_2;
  wire [0:0] muxN_1__in_data_3;
  wire [1:0] muxN_1__in_sel;
  wire [0:0] muxN_1__out;
  commonlib_muxn__N4__width1 muxN_1(
    .in_data_0(muxN_1__in_data_0),
    .in_data_1(muxN_1__in_data_1),
    .in_data_2(muxN_1__in_data_2),
    .in_data_3(muxN_1__in_data_3),
    .in_sel(muxN_1__in_sel),
    .out(muxN_1__out)
  );

  // Instancing generated Module: coreir.slice(hi:2, lo:0, width:3)
  wire [2:0] sel_slice0__in;
  wire [1:0] sel_slice0__out;
  coreir_slice #(.hi(2),.lo(0),.width(3)) sel_slice0(
    .in(sel_slice0__in),
    .out(sel_slice0__out)
  );

  // Instancing generated Module: coreir.slice(hi:2, lo:0, width:3)
  wire [2:0] sel_slice1__in;
  wire [1:0] sel_slice1__out;
  coreir_slice #(.hi(2),.lo(0),.width(3)) sel_slice1(
    .in(sel_slice1__in),
    .out(sel_slice1__out)
  );

  assign _join__in0[0:0] = muxN_0__out[0:0];

  assign _join__in1[0:0] = muxN_1__out[0:0];

  assign out[0:0] = _join__out[0:0];

  assign _join__sel = in_sel[2];

  assign muxN_0__in_data_0[0:0] = in_data_0[0:0];

  assign muxN_0__in_data_1[0:0] = in_data_1[0:0];

  assign muxN_0__in_data_2[0:0] = in_data_2[0:0];

  assign muxN_0__in_data_3[0:0] = in_data_3[0:0];

  assign muxN_0__in_sel[1:0] = sel_slice0__out[1:0];

  assign muxN_1__in_data_0[0:0] = in_data_4[0:0];

  assign muxN_1__in_data_1[0:0] = in_data_5[0:0];

  assign muxN_1__in_data_2[0:0] = in_data_6[0:0];

  assign muxN_1__in_data_3[0:0] = in_data_7[0:0];

  assign muxN_1__in_sel[1:0] = sel_slice1__out[1:0];

  assign sel_slice0__in[2:0] = in_sel[2:0];

  assign sel_slice1__in[2:0] = in_sel[2:0];


endmodule  // commonlib_muxn__N8__width1

// Generated from commonlib.muxn(N:1, width:32)
module commonlib_muxn__N1__width32 (
  input [31:0] in_data_0,
  input [0:0] in_sel,
  output [31:0] out
);


  wire  term_sel__in;
  corebit_term term_sel(
    .in(term_sel__in)
  );

  assign out[31:0] = in_data_0[31:0];

  assign term_sel__in = in_sel[0];


endmodule  // commonlib_muxn__N1__width32

// Generated from commonlib.muxn(N:3, width:32)
module commonlib_muxn__N3__width32 (
  input [31:0] in_data_0,
  input [31:0] in_data_1,
  input [31:0] in_data_2,
  input [1:0] in_sel,
  output [31:0] out
);


  // Instancing generated Module: coreir.mux(width:32)
  wire [31:0] _join__in0;
  wire [31:0] _join__in1;
  wire [31:0] _join__out;
  wire  _join__sel;
  coreir_mux #(.width(32)) _join(
    .in0(_join__in0),
    .in1(_join__in1),
    .out(_join__out),
    .sel(_join__sel)
  );

  // Instancing generated Module: commonlib.muxn(N:2, width:32)
  wire [31:0] muxN_0__in_data_0;
  wire [31:0] muxN_0__in_data_1;
  wire [0:0] muxN_0__in_sel;
  wire [31:0] muxN_0__out;
  commonlib_muxn__N2__width32 muxN_0(
    .in_data_0(muxN_0__in_data_0),
    .in_data_1(muxN_0__in_data_1),
    .in_sel(muxN_0__in_sel),
    .out(muxN_0__out)
  );

  // Instancing generated Module: commonlib.muxn(N:1, width:32)
  wire [31:0] muxN_1__in_data_0;
  wire [0:0] muxN_1__in_sel;
  wire [31:0] muxN_1__out;
  commonlib_muxn__N1__width32 muxN_1(
    .in_data_0(muxN_1__in_data_0),
    .in_sel(muxN_1__in_sel),
    .out(muxN_1__out)
  );

  // Instancing generated Module: coreir.slice(hi:1, lo:0, width:2)
  wire [1:0] sel_slice0__in;
  wire [0:0] sel_slice0__out;
  coreir_slice #(.hi(1),.lo(0),.width(2)) sel_slice0(
    .in(sel_slice0__in),
    .out(sel_slice0__out)
  );

  // Instancing generated Module: coreir.slice(hi:1, lo:0, width:2)
  wire [1:0] sel_slice1__in;
  wire [0:0] sel_slice1__out;
  coreir_slice #(.hi(1),.lo(0),.width(2)) sel_slice1(
    .in(sel_slice1__in),
    .out(sel_slice1__out)
  );

  assign _join__in0[31:0] = muxN_0__out[31:0];

  assign _join__in1[31:0] = muxN_1__out[31:0];

  assign out[31:0] = _join__out[31:0];

  assign _join__sel = in_sel[1];

  assign muxN_0__in_data_0[31:0] = in_data_0[31:0];

  assign muxN_0__in_data_1[31:0] = in_data_1[31:0];

  assign muxN_0__in_sel[0:0] = sel_slice0__out[0:0];

  assign muxN_1__in_data_0[31:0] = in_data_2[31:0];

  assign muxN_1__in_sel[0:0] = sel_slice1__out[0:0];

  assign sel_slice0__in[1:0] = in_sel[1:0];

  assign sel_slice1__in[1:0] = in_sel[1:0];


endmodule  // commonlib_muxn__N3__width32

// Generated from commonlib.muxn(N:7, width:32)
module commonlib_muxn__N7__width32 (
  input [31:0] in_data_0,
  input [31:0] in_data_1,
  input [31:0] in_data_2,
  input [31:0] in_data_3,
  input [31:0] in_data_4,
  input [31:0] in_data_5,
  input [31:0] in_data_6,
  input [2:0] in_sel,
  output [31:0] out
);


  // Instancing generated Module: coreir.mux(width:32)
  wire [31:0] _join__in0;
  wire [31:0] _join__in1;
  wire [31:0] _join__out;
  wire  _join__sel;
  coreir_mux #(.width(32)) _join(
    .in0(_join__in0),
    .in1(_join__in1),
    .out(_join__out),
    .sel(_join__sel)
  );

  // Instancing generated Module: commonlib.muxn(N:4, width:32)
  wire [31:0] muxN_0__in_data_0;
  wire [31:0] muxN_0__in_data_1;
  wire [31:0] muxN_0__in_data_2;
  wire [31:0] muxN_0__in_data_3;
  wire [1:0] muxN_0__in_sel;
  wire [31:0] muxN_0__out;
  commonlib_muxn__N4__width32 muxN_0(
    .in_data_0(muxN_0__in_data_0),
    .in_data_1(muxN_0__in_data_1),
    .in_data_2(muxN_0__in_data_2),
    .in_data_3(muxN_0__in_data_3),
    .in_sel(muxN_0__in_sel),
    .out(muxN_0__out)
  );

  // Instancing generated Module: commonlib.muxn(N:3, width:32)
  wire [31:0] muxN_1__in_data_0;
  wire [31:0] muxN_1__in_data_1;
  wire [31:0] muxN_1__in_data_2;
  wire [1:0] muxN_1__in_sel;
  wire [31:0] muxN_1__out;
  commonlib_muxn__N3__width32 muxN_1(
    .in_data_0(muxN_1__in_data_0),
    .in_data_1(muxN_1__in_data_1),
    .in_data_2(muxN_1__in_data_2),
    .in_sel(muxN_1__in_sel),
    .out(muxN_1__out)
  );

  // Instancing generated Module: coreir.slice(hi:2, lo:0, width:3)
  wire [2:0] sel_slice0__in;
  wire [1:0] sel_slice0__out;
  coreir_slice #(.hi(2),.lo(0),.width(3)) sel_slice0(
    .in(sel_slice0__in),
    .out(sel_slice0__out)
  );

  // Instancing generated Module: coreir.slice(hi:2, lo:0, width:3)
  wire [2:0] sel_slice1__in;
  wire [1:0] sel_slice1__out;
  coreir_slice #(.hi(2),.lo(0),.width(3)) sel_slice1(
    .in(sel_slice1__in),
    .out(sel_slice1__out)
  );

  assign _join__in0[31:0] = muxN_0__out[31:0];

  assign _join__in1[31:0] = muxN_1__out[31:0];

  assign out[31:0] = _join__out[31:0];

  assign _join__sel = in_sel[2];

  assign muxN_0__in_data_0[31:0] = in_data_0[31:0];

  assign muxN_0__in_data_1[31:0] = in_data_1[31:0];

  assign muxN_0__in_data_2[31:0] = in_data_2[31:0];

  assign muxN_0__in_data_3[31:0] = in_data_3[31:0];

  assign muxN_0__in_sel[1:0] = sel_slice0__out[1:0];

  assign muxN_1__in_data_0[31:0] = in_data_4[31:0];

  assign muxN_1__in_data_1[31:0] = in_data_5[31:0];

  assign muxN_1__in_data_2[31:0] = in_data_6[31:0];

  assign muxN_1__in_sel[1:0] = sel_slice1__out[1:0];

  assign sel_slice0__in[2:0] = in_sel[2:0];

  assign sel_slice1__in[2:0] = in_sel[2:0];


endmodule  // commonlib_muxn__N7__width32

// Generated from commonlib.muxn(N:16, width:32)
module commonlib_muxn__N16__width32 (
  input [31:0] in_data_0,
  input [31:0] in_data_1,
  input [31:0] in_data_10,
  input [31:0] in_data_11,
  input [31:0] in_data_12,
  input [31:0] in_data_13,
  input [31:0] in_data_14,
  input [31:0] in_data_15,
  input [31:0] in_data_2,
  input [31:0] in_data_3,
  input [31:0] in_data_4,
  input [31:0] in_data_5,
  input [31:0] in_data_6,
  input [31:0] in_data_7,
  input [31:0] in_data_8,
  input [31:0] in_data_9,
  input [3:0] in_sel,
  output [31:0] out
);


  // Instancing generated Module: coreir.mux(width:32)
  wire [31:0] _join__in0;
  wire [31:0] _join__in1;
  wire [31:0] _join__out;
  wire  _join__sel;
  coreir_mux #(.width(32)) _join(
    .in0(_join__in0),
    .in1(_join__in1),
    .out(_join__out),
    .sel(_join__sel)
  );

  // Instancing generated Module: commonlib.muxn(N:8, width:32)
  wire [31:0] muxN_0__in_data_0;
  wire [31:0] muxN_0__in_data_1;
  wire [31:0] muxN_0__in_data_2;
  wire [31:0] muxN_0__in_data_3;
  wire [31:0] muxN_0__in_data_4;
  wire [31:0] muxN_0__in_data_5;
  wire [31:0] muxN_0__in_data_6;
  wire [31:0] muxN_0__in_data_7;
  wire [2:0] muxN_0__in_sel;
  wire [31:0] muxN_0__out;
  commonlib_muxn__N8__width32 muxN_0(
    .in_data_0(muxN_0__in_data_0),
    .in_data_1(muxN_0__in_data_1),
    .in_data_2(muxN_0__in_data_2),
    .in_data_3(muxN_0__in_data_3),
    .in_data_4(muxN_0__in_data_4),
    .in_data_5(muxN_0__in_data_5),
    .in_data_6(muxN_0__in_data_6),
    .in_data_7(muxN_0__in_data_7),
    .in_sel(muxN_0__in_sel),
    .out(muxN_0__out)
  );

  // Instancing generated Module: commonlib.muxn(N:8, width:32)
  wire [31:0] muxN_1__in_data_0;
  wire [31:0] muxN_1__in_data_1;
  wire [31:0] muxN_1__in_data_2;
  wire [31:0] muxN_1__in_data_3;
  wire [31:0] muxN_1__in_data_4;
  wire [31:0] muxN_1__in_data_5;
  wire [31:0] muxN_1__in_data_6;
  wire [31:0] muxN_1__in_data_7;
  wire [2:0] muxN_1__in_sel;
  wire [31:0] muxN_1__out;
  commonlib_muxn__N8__width32 muxN_1(
    .in_data_0(muxN_1__in_data_0),
    .in_data_1(muxN_1__in_data_1),
    .in_data_2(muxN_1__in_data_2),
    .in_data_3(muxN_1__in_data_3),
    .in_data_4(muxN_1__in_data_4),
    .in_data_5(muxN_1__in_data_5),
    .in_data_6(muxN_1__in_data_6),
    .in_data_7(muxN_1__in_data_7),
    .in_sel(muxN_1__in_sel),
    .out(muxN_1__out)
  );

  // Instancing generated Module: coreir.slice(hi:3, lo:0, width:4)
  wire [3:0] sel_slice0__in;
  wire [2:0] sel_slice0__out;
  coreir_slice #(.hi(3),.lo(0),.width(4)) sel_slice0(
    .in(sel_slice0__in),
    .out(sel_slice0__out)
  );

  // Instancing generated Module: coreir.slice(hi:3, lo:0, width:4)
  wire [3:0] sel_slice1__in;
  wire [2:0] sel_slice1__out;
  coreir_slice #(.hi(3),.lo(0),.width(4)) sel_slice1(
    .in(sel_slice1__in),
    .out(sel_slice1__out)
  );

  assign _join__in0[31:0] = muxN_0__out[31:0];

  assign _join__in1[31:0] = muxN_1__out[31:0];

  assign out[31:0] = _join__out[31:0];

  assign _join__sel = in_sel[3];

  assign muxN_0__in_data_0[31:0] = in_data_0[31:0];

  assign muxN_0__in_data_1[31:0] = in_data_1[31:0];

  assign muxN_0__in_data_2[31:0] = in_data_2[31:0];

  assign muxN_0__in_data_3[31:0] = in_data_3[31:0];

  assign muxN_0__in_data_4[31:0] = in_data_4[31:0];

  assign muxN_0__in_data_5[31:0] = in_data_5[31:0];

  assign muxN_0__in_data_6[31:0] = in_data_6[31:0];

  assign muxN_0__in_data_7[31:0] = in_data_7[31:0];

  assign muxN_0__in_sel[2:0] = sel_slice0__out[2:0];

  assign muxN_1__in_data_0[31:0] = in_data_8[31:0];

  assign muxN_1__in_data_1[31:0] = in_data_9[31:0];

  assign muxN_1__in_data_2[31:0] = in_data_10[31:0];

  assign muxN_1__in_data_3[31:0] = in_data_11[31:0];

  assign muxN_1__in_data_4[31:0] = in_data_12[31:0];

  assign muxN_1__in_data_5[31:0] = in_data_13[31:0];

  assign muxN_1__in_data_6[31:0] = in_data_14[31:0];

  assign muxN_1__in_data_7[31:0] = in_data_15[31:0];

  assign muxN_1__in_sel[2:0] = sel_slice1__out[2:0];

  assign sel_slice0__in[3:0] = in_sel[3:0];

  assign sel_slice1__in[3:0] = in_sel[3:0];


endmodule  // commonlib_muxn__N16__width32

// Generated from commonlib.muxn(N:32, width:32)
module commonlib_muxn__N32__width32 (
  input [31:0] in_data_0,
  input [31:0] in_data_1,
  input [31:0] in_data_10,
  input [31:0] in_data_11,
  input [31:0] in_data_12,
  input [31:0] in_data_13,
  input [31:0] in_data_14,
  input [31:0] in_data_15,
  input [31:0] in_data_16,
  input [31:0] in_data_17,
  input [31:0] in_data_18,
  input [31:0] in_data_19,
  input [31:0] in_data_2,
  input [31:0] in_data_20,
  input [31:0] in_data_21,
  input [31:0] in_data_22,
  input [31:0] in_data_23,
  input [31:0] in_data_24,
  input [31:0] in_data_25,
  input [31:0] in_data_26,
  input [31:0] in_data_27,
  input [31:0] in_data_28,
  input [31:0] in_data_29,
  input [31:0] in_data_3,
  input [31:0] in_data_30,
  input [31:0] in_data_31,
  input [31:0] in_data_4,
  input [31:0] in_data_5,
  input [31:0] in_data_6,
  input [31:0] in_data_7,
  input [31:0] in_data_8,
  input [31:0] in_data_9,
  input [4:0] in_sel,
  output [31:0] out
);


  // Instancing generated Module: coreir.mux(width:32)
  wire [31:0] _join__in0;
  wire [31:0] _join__in1;
  wire [31:0] _join__out;
  wire  _join__sel;
  coreir_mux #(.width(32)) _join(
    .in0(_join__in0),
    .in1(_join__in1),
    .out(_join__out),
    .sel(_join__sel)
  );

  // Instancing generated Module: commonlib.muxn(N:16, width:32)
  wire [31:0] muxN_0__in_data_0;
  wire [31:0] muxN_0__in_data_1;
  wire [31:0] muxN_0__in_data_10;
  wire [31:0] muxN_0__in_data_11;
  wire [31:0] muxN_0__in_data_12;
  wire [31:0] muxN_0__in_data_13;
  wire [31:0] muxN_0__in_data_14;
  wire [31:0] muxN_0__in_data_15;
  wire [31:0] muxN_0__in_data_2;
  wire [31:0] muxN_0__in_data_3;
  wire [31:0] muxN_0__in_data_4;
  wire [31:0] muxN_0__in_data_5;
  wire [31:0] muxN_0__in_data_6;
  wire [31:0] muxN_0__in_data_7;
  wire [31:0] muxN_0__in_data_8;
  wire [31:0] muxN_0__in_data_9;
  wire [3:0] muxN_0__in_sel;
  wire [31:0] muxN_0__out;
  commonlib_muxn__N16__width32 muxN_0(
    .in_data_0(muxN_0__in_data_0),
    .in_data_1(muxN_0__in_data_1),
    .in_data_10(muxN_0__in_data_10),
    .in_data_11(muxN_0__in_data_11),
    .in_data_12(muxN_0__in_data_12),
    .in_data_13(muxN_0__in_data_13),
    .in_data_14(muxN_0__in_data_14),
    .in_data_15(muxN_0__in_data_15),
    .in_data_2(muxN_0__in_data_2),
    .in_data_3(muxN_0__in_data_3),
    .in_data_4(muxN_0__in_data_4),
    .in_data_5(muxN_0__in_data_5),
    .in_data_6(muxN_0__in_data_6),
    .in_data_7(muxN_0__in_data_7),
    .in_data_8(muxN_0__in_data_8),
    .in_data_9(muxN_0__in_data_9),
    .in_sel(muxN_0__in_sel),
    .out(muxN_0__out)
  );

  // Instancing generated Module: commonlib.muxn(N:16, width:32)
  wire [31:0] muxN_1__in_data_0;
  wire [31:0] muxN_1__in_data_1;
  wire [31:0] muxN_1__in_data_10;
  wire [31:0] muxN_1__in_data_11;
  wire [31:0] muxN_1__in_data_12;
  wire [31:0] muxN_1__in_data_13;
  wire [31:0] muxN_1__in_data_14;
  wire [31:0] muxN_1__in_data_15;
  wire [31:0] muxN_1__in_data_2;
  wire [31:0] muxN_1__in_data_3;
  wire [31:0] muxN_1__in_data_4;
  wire [31:0] muxN_1__in_data_5;
  wire [31:0] muxN_1__in_data_6;
  wire [31:0] muxN_1__in_data_7;
  wire [31:0] muxN_1__in_data_8;
  wire [31:0] muxN_1__in_data_9;
  wire [3:0] muxN_1__in_sel;
  wire [31:0] muxN_1__out;
  commonlib_muxn__N16__width32 muxN_1(
    .in_data_0(muxN_1__in_data_0),
    .in_data_1(muxN_1__in_data_1),
    .in_data_10(muxN_1__in_data_10),
    .in_data_11(muxN_1__in_data_11),
    .in_data_12(muxN_1__in_data_12),
    .in_data_13(muxN_1__in_data_13),
    .in_data_14(muxN_1__in_data_14),
    .in_data_15(muxN_1__in_data_15),
    .in_data_2(muxN_1__in_data_2),
    .in_data_3(muxN_1__in_data_3),
    .in_data_4(muxN_1__in_data_4),
    .in_data_5(muxN_1__in_data_5),
    .in_data_6(muxN_1__in_data_6),
    .in_data_7(muxN_1__in_data_7),
    .in_data_8(muxN_1__in_data_8),
    .in_data_9(muxN_1__in_data_9),
    .in_sel(muxN_1__in_sel),
    .out(muxN_1__out)
  );

  // Instancing generated Module: coreir.slice(hi:4, lo:0, width:5)
  wire [4:0] sel_slice0__in;
  wire [3:0] sel_slice0__out;
  coreir_slice #(.hi(4),.lo(0),.width(5)) sel_slice0(
    .in(sel_slice0__in),
    .out(sel_slice0__out)
  );

  // Instancing generated Module: coreir.slice(hi:4, lo:0, width:5)
  wire [4:0] sel_slice1__in;
  wire [3:0] sel_slice1__out;
  coreir_slice #(.hi(4),.lo(0),.width(5)) sel_slice1(
    .in(sel_slice1__in),
    .out(sel_slice1__out)
  );

  assign _join__in0[31:0] = muxN_0__out[31:0];

  assign _join__in1[31:0] = muxN_1__out[31:0];

  assign out[31:0] = _join__out[31:0];

  assign _join__sel = in_sel[4];

  assign muxN_0__in_data_0[31:0] = in_data_0[31:0];

  assign muxN_0__in_data_1[31:0] = in_data_1[31:0];

  assign muxN_0__in_data_10[31:0] = in_data_10[31:0];

  assign muxN_0__in_data_11[31:0] = in_data_11[31:0];

  assign muxN_0__in_data_12[31:0] = in_data_12[31:0];

  assign muxN_0__in_data_13[31:0] = in_data_13[31:0];

  assign muxN_0__in_data_14[31:0] = in_data_14[31:0];

  assign muxN_0__in_data_15[31:0] = in_data_15[31:0];

  assign muxN_0__in_data_2[31:0] = in_data_2[31:0];

  assign muxN_0__in_data_3[31:0] = in_data_3[31:0];

  assign muxN_0__in_data_4[31:0] = in_data_4[31:0];

  assign muxN_0__in_data_5[31:0] = in_data_5[31:0];

  assign muxN_0__in_data_6[31:0] = in_data_6[31:0];

  assign muxN_0__in_data_7[31:0] = in_data_7[31:0];

  assign muxN_0__in_data_8[31:0] = in_data_8[31:0];

  assign muxN_0__in_data_9[31:0] = in_data_9[31:0];

  assign muxN_0__in_sel[3:0] = sel_slice0__out[3:0];

  assign muxN_1__in_data_0[31:0] = in_data_16[31:0];

  assign muxN_1__in_data_1[31:0] = in_data_17[31:0];

  assign muxN_1__in_data_10[31:0] = in_data_26[31:0];

  assign muxN_1__in_data_11[31:0] = in_data_27[31:0];

  assign muxN_1__in_data_12[31:0] = in_data_28[31:0];

  assign muxN_1__in_data_13[31:0] = in_data_29[31:0];

  assign muxN_1__in_data_14[31:0] = in_data_30[31:0];

  assign muxN_1__in_data_15[31:0] = in_data_31[31:0];

  assign muxN_1__in_data_2[31:0] = in_data_18[31:0];

  assign muxN_1__in_data_3[31:0] = in_data_19[31:0];

  assign muxN_1__in_data_4[31:0] = in_data_20[31:0];

  assign muxN_1__in_data_5[31:0] = in_data_21[31:0];

  assign muxN_1__in_data_6[31:0] = in_data_22[31:0];

  assign muxN_1__in_data_7[31:0] = in_data_23[31:0];

  assign muxN_1__in_data_8[31:0] = in_data_24[31:0];

  assign muxN_1__in_data_9[31:0] = in_data_25[31:0];

  assign muxN_1__in_sel[3:0] = sel_slice1__out[3:0];

  assign sel_slice0__in[4:0] = in_sel[4:0];

  assign sel_slice1__in[4:0] = in_sel[4:0];


endmodule  // commonlib_muxn__N32__width32

// Generated from commonlib.muxn(N:64, width:32)
module commonlib_muxn__N64__width32 (
  input [31:0] in_data_0,
  input [31:0] in_data_1,
  input [31:0] in_data_10,
  input [31:0] in_data_11,
  input [31:0] in_data_12,
  input [31:0] in_data_13,
  input [31:0] in_data_14,
  input [31:0] in_data_15,
  input [31:0] in_data_16,
  input [31:0] in_data_17,
  input [31:0] in_data_18,
  input [31:0] in_data_19,
  input [31:0] in_data_2,
  input [31:0] in_data_20,
  input [31:0] in_data_21,
  input [31:0] in_data_22,
  input [31:0] in_data_23,
  input [31:0] in_data_24,
  input [31:0] in_data_25,
  input [31:0] in_data_26,
  input [31:0] in_data_27,
  input [31:0] in_data_28,
  input [31:0] in_data_29,
  input [31:0] in_data_3,
  input [31:0] in_data_30,
  input [31:0] in_data_31,
  input [31:0] in_data_32,
  input [31:0] in_data_33,
  input [31:0] in_data_34,
  input [31:0] in_data_35,
  input [31:0] in_data_36,
  input [31:0] in_data_37,
  input [31:0] in_data_38,
  input [31:0] in_data_39,
  input [31:0] in_data_4,
  input [31:0] in_data_40,
  input [31:0] in_data_41,
  input [31:0] in_data_42,
  input [31:0] in_data_43,
  input [31:0] in_data_44,
  input [31:0] in_data_45,
  input [31:0] in_data_46,
  input [31:0] in_data_47,
  input [31:0] in_data_48,
  input [31:0] in_data_49,
  input [31:0] in_data_5,
  input [31:0] in_data_50,
  input [31:0] in_data_51,
  input [31:0] in_data_52,
  input [31:0] in_data_53,
  input [31:0] in_data_54,
  input [31:0] in_data_55,
  input [31:0] in_data_56,
  input [31:0] in_data_57,
  input [31:0] in_data_58,
  input [31:0] in_data_59,
  input [31:0] in_data_6,
  input [31:0] in_data_60,
  input [31:0] in_data_61,
  input [31:0] in_data_62,
  input [31:0] in_data_63,
  input [31:0] in_data_7,
  input [31:0] in_data_8,
  input [31:0] in_data_9,
  input [5:0] in_sel,
  output [31:0] out
);


  // Instancing generated Module: coreir.mux(width:32)
  wire [31:0] _join__in0;
  wire [31:0] _join__in1;
  wire [31:0] _join__out;
  wire  _join__sel;
  coreir_mux #(.width(32)) _join(
    .in0(_join__in0),
    .in1(_join__in1),
    .out(_join__out),
    .sel(_join__sel)
  );

  // Instancing generated Module: commonlib.muxn(N:32, width:32)
  wire [31:0] muxN_0__in_data_0;
  wire [31:0] muxN_0__in_data_1;
  wire [31:0] muxN_0__in_data_10;
  wire [31:0] muxN_0__in_data_11;
  wire [31:0] muxN_0__in_data_12;
  wire [31:0] muxN_0__in_data_13;
  wire [31:0] muxN_0__in_data_14;
  wire [31:0] muxN_0__in_data_15;
  wire [31:0] muxN_0__in_data_16;
  wire [31:0] muxN_0__in_data_17;
  wire [31:0] muxN_0__in_data_18;
  wire [31:0] muxN_0__in_data_19;
  wire [31:0] muxN_0__in_data_2;
  wire [31:0] muxN_0__in_data_20;
  wire [31:0] muxN_0__in_data_21;
  wire [31:0] muxN_0__in_data_22;
  wire [31:0] muxN_0__in_data_23;
  wire [31:0] muxN_0__in_data_24;
  wire [31:0] muxN_0__in_data_25;
  wire [31:0] muxN_0__in_data_26;
  wire [31:0] muxN_0__in_data_27;
  wire [31:0] muxN_0__in_data_28;
  wire [31:0] muxN_0__in_data_29;
  wire [31:0] muxN_0__in_data_3;
  wire [31:0] muxN_0__in_data_30;
  wire [31:0] muxN_0__in_data_31;
  wire [31:0] muxN_0__in_data_4;
  wire [31:0] muxN_0__in_data_5;
  wire [31:0] muxN_0__in_data_6;
  wire [31:0] muxN_0__in_data_7;
  wire [31:0] muxN_0__in_data_8;
  wire [31:0] muxN_0__in_data_9;
  wire [4:0] muxN_0__in_sel;
  wire [31:0] muxN_0__out;
  commonlib_muxn__N32__width32 muxN_0(
    .in_data_0(muxN_0__in_data_0),
    .in_data_1(muxN_0__in_data_1),
    .in_data_10(muxN_0__in_data_10),
    .in_data_11(muxN_0__in_data_11),
    .in_data_12(muxN_0__in_data_12),
    .in_data_13(muxN_0__in_data_13),
    .in_data_14(muxN_0__in_data_14),
    .in_data_15(muxN_0__in_data_15),
    .in_data_16(muxN_0__in_data_16),
    .in_data_17(muxN_0__in_data_17),
    .in_data_18(muxN_0__in_data_18),
    .in_data_19(muxN_0__in_data_19),
    .in_data_2(muxN_0__in_data_2),
    .in_data_20(muxN_0__in_data_20),
    .in_data_21(muxN_0__in_data_21),
    .in_data_22(muxN_0__in_data_22),
    .in_data_23(muxN_0__in_data_23),
    .in_data_24(muxN_0__in_data_24),
    .in_data_25(muxN_0__in_data_25),
    .in_data_26(muxN_0__in_data_26),
    .in_data_27(muxN_0__in_data_27),
    .in_data_28(muxN_0__in_data_28),
    .in_data_29(muxN_0__in_data_29),
    .in_data_3(muxN_0__in_data_3),
    .in_data_30(muxN_0__in_data_30),
    .in_data_31(muxN_0__in_data_31),
    .in_data_4(muxN_0__in_data_4),
    .in_data_5(muxN_0__in_data_5),
    .in_data_6(muxN_0__in_data_6),
    .in_data_7(muxN_0__in_data_7),
    .in_data_8(muxN_0__in_data_8),
    .in_data_9(muxN_0__in_data_9),
    .in_sel(muxN_0__in_sel),
    .out(muxN_0__out)
  );

  // Instancing generated Module: commonlib.muxn(N:32, width:32)
  wire [31:0] muxN_1__in_data_0;
  wire [31:0] muxN_1__in_data_1;
  wire [31:0] muxN_1__in_data_10;
  wire [31:0] muxN_1__in_data_11;
  wire [31:0] muxN_1__in_data_12;
  wire [31:0] muxN_1__in_data_13;
  wire [31:0] muxN_1__in_data_14;
  wire [31:0] muxN_1__in_data_15;
  wire [31:0] muxN_1__in_data_16;
  wire [31:0] muxN_1__in_data_17;
  wire [31:0] muxN_1__in_data_18;
  wire [31:0] muxN_1__in_data_19;
  wire [31:0] muxN_1__in_data_2;
  wire [31:0] muxN_1__in_data_20;
  wire [31:0] muxN_1__in_data_21;
  wire [31:0] muxN_1__in_data_22;
  wire [31:0] muxN_1__in_data_23;
  wire [31:0] muxN_1__in_data_24;
  wire [31:0] muxN_1__in_data_25;
  wire [31:0] muxN_1__in_data_26;
  wire [31:0] muxN_1__in_data_27;
  wire [31:0] muxN_1__in_data_28;
  wire [31:0] muxN_1__in_data_29;
  wire [31:0] muxN_1__in_data_3;
  wire [31:0] muxN_1__in_data_30;
  wire [31:0] muxN_1__in_data_31;
  wire [31:0] muxN_1__in_data_4;
  wire [31:0] muxN_1__in_data_5;
  wire [31:0] muxN_1__in_data_6;
  wire [31:0] muxN_1__in_data_7;
  wire [31:0] muxN_1__in_data_8;
  wire [31:0] muxN_1__in_data_9;
  wire [4:0] muxN_1__in_sel;
  wire [31:0] muxN_1__out;
  commonlib_muxn__N32__width32 muxN_1(
    .in_data_0(muxN_1__in_data_0),
    .in_data_1(muxN_1__in_data_1),
    .in_data_10(muxN_1__in_data_10),
    .in_data_11(muxN_1__in_data_11),
    .in_data_12(muxN_1__in_data_12),
    .in_data_13(muxN_1__in_data_13),
    .in_data_14(muxN_1__in_data_14),
    .in_data_15(muxN_1__in_data_15),
    .in_data_16(muxN_1__in_data_16),
    .in_data_17(muxN_1__in_data_17),
    .in_data_18(muxN_1__in_data_18),
    .in_data_19(muxN_1__in_data_19),
    .in_data_2(muxN_1__in_data_2),
    .in_data_20(muxN_1__in_data_20),
    .in_data_21(muxN_1__in_data_21),
    .in_data_22(muxN_1__in_data_22),
    .in_data_23(muxN_1__in_data_23),
    .in_data_24(muxN_1__in_data_24),
    .in_data_25(muxN_1__in_data_25),
    .in_data_26(muxN_1__in_data_26),
    .in_data_27(muxN_1__in_data_27),
    .in_data_28(muxN_1__in_data_28),
    .in_data_29(muxN_1__in_data_29),
    .in_data_3(muxN_1__in_data_3),
    .in_data_30(muxN_1__in_data_30),
    .in_data_31(muxN_1__in_data_31),
    .in_data_4(muxN_1__in_data_4),
    .in_data_5(muxN_1__in_data_5),
    .in_data_6(muxN_1__in_data_6),
    .in_data_7(muxN_1__in_data_7),
    .in_data_8(muxN_1__in_data_8),
    .in_data_9(muxN_1__in_data_9),
    .in_sel(muxN_1__in_sel),
    .out(muxN_1__out)
  );

  // Instancing generated Module: coreir.slice(hi:5, lo:0, width:6)
  wire [5:0] sel_slice0__in;
  wire [4:0] sel_slice0__out;
  coreir_slice #(.hi(5),.lo(0),.width(6)) sel_slice0(
    .in(sel_slice0__in),
    .out(sel_slice0__out)
  );

  // Instancing generated Module: coreir.slice(hi:5, lo:0, width:6)
  wire [5:0] sel_slice1__in;
  wire [4:0] sel_slice1__out;
  coreir_slice #(.hi(5),.lo(0),.width(6)) sel_slice1(
    .in(sel_slice1__in),
    .out(sel_slice1__out)
  );

  assign _join__in0[31:0] = muxN_0__out[31:0];

  assign _join__in1[31:0] = muxN_1__out[31:0];

  assign out[31:0] = _join__out[31:0];

  assign _join__sel = in_sel[5];

  assign muxN_0__in_data_0[31:0] = in_data_0[31:0];

  assign muxN_0__in_data_1[31:0] = in_data_1[31:0];

  assign muxN_0__in_data_10[31:0] = in_data_10[31:0];

  assign muxN_0__in_data_11[31:0] = in_data_11[31:0];

  assign muxN_0__in_data_12[31:0] = in_data_12[31:0];

  assign muxN_0__in_data_13[31:0] = in_data_13[31:0];

  assign muxN_0__in_data_14[31:0] = in_data_14[31:0];

  assign muxN_0__in_data_15[31:0] = in_data_15[31:0];

  assign muxN_0__in_data_16[31:0] = in_data_16[31:0];

  assign muxN_0__in_data_17[31:0] = in_data_17[31:0];

  assign muxN_0__in_data_18[31:0] = in_data_18[31:0];

  assign muxN_0__in_data_19[31:0] = in_data_19[31:0];

  assign muxN_0__in_data_2[31:0] = in_data_2[31:0];

  assign muxN_0__in_data_20[31:0] = in_data_20[31:0];

  assign muxN_0__in_data_21[31:0] = in_data_21[31:0];

  assign muxN_0__in_data_22[31:0] = in_data_22[31:0];

  assign muxN_0__in_data_23[31:0] = in_data_23[31:0];

  assign muxN_0__in_data_24[31:0] = in_data_24[31:0];

  assign muxN_0__in_data_25[31:0] = in_data_25[31:0];

  assign muxN_0__in_data_26[31:0] = in_data_26[31:0];

  assign muxN_0__in_data_27[31:0] = in_data_27[31:0];

  assign muxN_0__in_data_28[31:0] = in_data_28[31:0];

  assign muxN_0__in_data_29[31:0] = in_data_29[31:0];

  assign muxN_0__in_data_3[31:0] = in_data_3[31:0];

  assign muxN_0__in_data_30[31:0] = in_data_30[31:0];

  assign muxN_0__in_data_31[31:0] = in_data_31[31:0];

  assign muxN_0__in_data_4[31:0] = in_data_4[31:0];

  assign muxN_0__in_data_5[31:0] = in_data_5[31:0];

  assign muxN_0__in_data_6[31:0] = in_data_6[31:0];

  assign muxN_0__in_data_7[31:0] = in_data_7[31:0];

  assign muxN_0__in_data_8[31:0] = in_data_8[31:0];

  assign muxN_0__in_data_9[31:0] = in_data_9[31:0];

  assign muxN_0__in_sel[4:0] = sel_slice0__out[4:0];

  assign muxN_1__in_data_0[31:0] = in_data_32[31:0];

  assign muxN_1__in_data_1[31:0] = in_data_33[31:0];

  assign muxN_1__in_data_10[31:0] = in_data_42[31:0];

  assign muxN_1__in_data_11[31:0] = in_data_43[31:0];

  assign muxN_1__in_data_12[31:0] = in_data_44[31:0];

  assign muxN_1__in_data_13[31:0] = in_data_45[31:0];

  assign muxN_1__in_data_14[31:0] = in_data_46[31:0];

  assign muxN_1__in_data_15[31:0] = in_data_47[31:0];

  assign muxN_1__in_data_16[31:0] = in_data_48[31:0];

  assign muxN_1__in_data_17[31:0] = in_data_49[31:0];

  assign muxN_1__in_data_18[31:0] = in_data_50[31:0];

  assign muxN_1__in_data_19[31:0] = in_data_51[31:0];

  assign muxN_1__in_data_2[31:0] = in_data_34[31:0];

  assign muxN_1__in_data_20[31:0] = in_data_52[31:0];

  assign muxN_1__in_data_21[31:0] = in_data_53[31:0];

  assign muxN_1__in_data_22[31:0] = in_data_54[31:0];

  assign muxN_1__in_data_23[31:0] = in_data_55[31:0];

  assign muxN_1__in_data_24[31:0] = in_data_56[31:0];

  assign muxN_1__in_data_25[31:0] = in_data_57[31:0];

  assign muxN_1__in_data_26[31:0] = in_data_58[31:0];

  assign muxN_1__in_data_27[31:0] = in_data_59[31:0];

  assign muxN_1__in_data_28[31:0] = in_data_60[31:0];

  assign muxN_1__in_data_29[31:0] = in_data_61[31:0];

  assign muxN_1__in_data_3[31:0] = in_data_35[31:0];

  assign muxN_1__in_data_30[31:0] = in_data_62[31:0];

  assign muxN_1__in_data_31[31:0] = in_data_63[31:0];

  assign muxN_1__in_data_4[31:0] = in_data_36[31:0];

  assign muxN_1__in_data_5[31:0] = in_data_37[31:0];

  assign muxN_1__in_data_6[31:0] = in_data_38[31:0];

  assign muxN_1__in_data_7[31:0] = in_data_39[31:0];

  assign muxN_1__in_data_8[31:0] = in_data_40[31:0];

  assign muxN_1__in_data_9[31:0] = in_data_41[31:0];

  assign muxN_1__in_sel[4:0] = sel_slice1__out[4:0];

  assign sel_slice0__in[5:0] = in_sel[5:0];

  assign sel_slice1__in[5:0] = in_sel[5:0];


endmodule  // commonlib_muxn__N64__width32

// Generated from commonlib.muxn(N:80, width:32)
module commonlib_muxn__N80__width32 (
  input [31:0] in_data_0,
  input [31:0] in_data_1,
  input [31:0] in_data_10,
  input [31:0] in_data_11,
  input [31:0] in_data_12,
  input [31:0] in_data_13,
  input [31:0] in_data_14,
  input [31:0] in_data_15,
  input [31:0] in_data_16,
  input [31:0] in_data_17,
  input [31:0] in_data_18,
  input [31:0] in_data_19,
  input [31:0] in_data_2,
  input [31:0] in_data_20,
  input [31:0] in_data_21,
  input [31:0] in_data_22,
  input [31:0] in_data_23,
  input [31:0] in_data_24,
  input [31:0] in_data_25,
  input [31:0] in_data_26,
  input [31:0] in_data_27,
  input [31:0] in_data_28,
  input [31:0] in_data_29,
  input [31:0] in_data_3,
  input [31:0] in_data_30,
  input [31:0] in_data_31,
  input [31:0] in_data_32,
  input [31:0] in_data_33,
  input [31:0] in_data_34,
  input [31:0] in_data_35,
  input [31:0] in_data_36,
  input [31:0] in_data_37,
  input [31:0] in_data_38,
  input [31:0] in_data_39,
  input [31:0] in_data_4,
  input [31:0] in_data_40,
  input [31:0] in_data_41,
  input [31:0] in_data_42,
  input [31:0] in_data_43,
  input [31:0] in_data_44,
  input [31:0] in_data_45,
  input [31:0] in_data_46,
  input [31:0] in_data_47,
  input [31:0] in_data_48,
  input [31:0] in_data_49,
  input [31:0] in_data_5,
  input [31:0] in_data_50,
  input [31:0] in_data_51,
  input [31:0] in_data_52,
  input [31:0] in_data_53,
  input [31:0] in_data_54,
  input [31:0] in_data_55,
  input [31:0] in_data_56,
  input [31:0] in_data_57,
  input [31:0] in_data_58,
  input [31:0] in_data_59,
  input [31:0] in_data_6,
  input [31:0] in_data_60,
  input [31:0] in_data_61,
  input [31:0] in_data_62,
  input [31:0] in_data_63,
  input [31:0] in_data_64,
  input [31:0] in_data_65,
  input [31:0] in_data_66,
  input [31:0] in_data_67,
  input [31:0] in_data_68,
  input [31:0] in_data_69,
  input [31:0] in_data_7,
  input [31:0] in_data_70,
  input [31:0] in_data_71,
  input [31:0] in_data_72,
  input [31:0] in_data_73,
  input [31:0] in_data_74,
  input [31:0] in_data_75,
  input [31:0] in_data_76,
  input [31:0] in_data_77,
  input [31:0] in_data_78,
  input [31:0] in_data_79,
  input [31:0] in_data_8,
  input [31:0] in_data_9,
  input [6:0] in_sel,
  output [31:0] out
);


  // Instancing generated Module: coreir.mux(width:32)
  wire [31:0] _join__in0;
  wire [31:0] _join__in1;
  wire [31:0] _join__out;
  wire  _join__sel;
  coreir_mux #(.width(32)) _join(
    .in0(_join__in0),
    .in1(_join__in1),
    .out(_join__out),
    .sel(_join__sel)
  );

  // Instancing generated Module: commonlib.muxn(N:64, width:32)
  wire [31:0] muxN_0__in_data_0;
  wire [31:0] muxN_0__in_data_1;
  wire [31:0] muxN_0__in_data_10;
  wire [31:0] muxN_0__in_data_11;
  wire [31:0] muxN_0__in_data_12;
  wire [31:0] muxN_0__in_data_13;
  wire [31:0] muxN_0__in_data_14;
  wire [31:0] muxN_0__in_data_15;
  wire [31:0] muxN_0__in_data_16;
  wire [31:0] muxN_0__in_data_17;
  wire [31:0] muxN_0__in_data_18;
  wire [31:0] muxN_0__in_data_19;
  wire [31:0] muxN_0__in_data_2;
  wire [31:0] muxN_0__in_data_20;
  wire [31:0] muxN_0__in_data_21;
  wire [31:0] muxN_0__in_data_22;
  wire [31:0] muxN_0__in_data_23;
  wire [31:0] muxN_0__in_data_24;
  wire [31:0] muxN_0__in_data_25;
  wire [31:0] muxN_0__in_data_26;
  wire [31:0] muxN_0__in_data_27;
  wire [31:0] muxN_0__in_data_28;
  wire [31:0] muxN_0__in_data_29;
  wire [31:0] muxN_0__in_data_3;
  wire [31:0] muxN_0__in_data_30;
  wire [31:0] muxN_0__in_data_31;
  wire [31:0] muxN_0__in_data_32;
  wire [31:0] muxN_0__in_data_33;
  wire [31:0] muxN_0__in_data_34;
  wire [31:0] muxN_0__in_data_35;
  wire [31:0] muxN_0__in_data_36;
  wire [31:0] muxN_0__in_data_37;
  wire [31:0] muxN_0__in_data_38;
  wire [31:0] muxN_0__in_data_39;
  wire [31:0] muxN_0__in_data_4;
  wire [31:0] muxN_0__in_data_40;
  wire [31:0] muxN_0__in_data_41;
  wire [31:0] muxN_0__in_data_42;
  wire [31:0] muxN_0__in_data_43;
  wire [31:0] muxN_0__in_data_44;
  wire [31:0] muxN_0__in_data_45;
  wire [31:0] muxN_0__in_data_46;
  wire [31:0] muxN_0__in_data_47;
  wire [31:0] muxN_0__in_data_48;
  wire [31:0] muxN_0__in_data_49;
  wire [31:0] muxN_0__in_data_5;
  wire [31:0] muxN_0__in_data_50;
  wire [31:0] muxN_0__in_data_51;
  wire [31:0] muxN_0__in_data_52;
  wire [31:0] muxN_0__in_data_53;
  wire [31:0] muxN_0__in_data_54;
  wire [31:0] muxN_0__in_data_55;
  wire [31:0] muxN_0__in_data_56;
  wire [31:0] muxN_0__in_data_57;
  wire [31:0] muxN_0__in_data_58;
  wire [31:0] muxN_0__in_data_59;
  wire [31:0] muxN_0__in_data_6;
  wire [31:0] muxN_0__in_data_60;
  wire [31:0] muxN_0__in_data_61;
  wire [31:0] muxN_0__in_data_62;
  wire [31:0] muxN_0__in_data_63;
  wire [31:0] muxN_0__in_data_7;
  wire [31:0] muxN_0__in_data_8;
  wire [31:0] muxN_0__in_data_9;
  wire [5:0] muxN_0__in_sel;
  wire [31:0] muxN_0__out;
  commonlib_muxn__N64__width32 muxN_0(
    .in_data_0(muxN_0__in_data_0),
    .in_data_1(muxN_0__in_data_1),
    .in_data_10(muxN_0__in_data_10),
    .in_data_11(muxN_0__in_data_11),
    .in_data_12(muxN_0__in_data_12),
    .in_data_13(muxN_0__in_data_13),
    .in_data_14(muxN_0__in_data_14),
    .in_data_15(muxN_0__in_data_15),
    .in_data_16(muxN_0__in_data_16),
    .in_data_17(muxN_0__in_data_17),
    .in_data_18(muxN_0__in_data_18),
    .in_data_19(muxN_0__in_data_19),
    .in_data_2(muxN_0__in_data_2),
    .in_data_20(muxN_0__in_data_20),
    .in_data_21(muxN_0__in_data_21),
    .in_data_22(muxN_0__in_data_22),
    .in_data_23(muxN_0__in_data_23),
    .in_data_24(muxN_0__in_data_24),
    .in_data_25(muxN_0__in_data_25),
    .in_data_26(muxN_0__in_data_26),
    .in_data_27(muxN_0__in_data_27),
    .in_data_28(muxN_0__in_data_28),
    .in_data_29(muxN_0__in_data_29),
    .in_data_3(muxN_0__in_data_3),
    .in_data_30(muxN_0__in_data_30),
    .in_data_31(muxN_0__in_data_31),
    .in_data_32(muxN_0__in_data_32),
    .in_data_33(muxN_0__in_data_33),
    .in_data_34(muxN_0__in_data_34),
    .in_data_35(muxN_0__in_data_35),
    .in_data_36(muxN_0__in_data_36),
    .in_data_37(muxN_0__in_data_37),
    .in_data_38(muxN_0__in_data_38),
    .in_data_39(muxN_0__in_data_39),
    .in_data_4(muxN_0__in_data_4),
    .in_data_40(muxN_0__in_data_40),
    .in_data_41(muxN_0__in_data_41),
    .in_data_42(muxN_0__in_data_42),
    .in_data_43(muxN_0__in_data_43),
    .in_data_44(muxN_0__in_data_44),
    .in_data_45(muxN_0__in_data_45),
    .in_data_46(muxN_0__in_data_46),
    .in_data_47(muxN_0__in_data_47),
    .in_data_48(muxN_0__in_data_48),
    .in_data_49(muxN_0__in_data_49),
    .in_data_5(muxN_0__in_data_5),
    .in_data_50(muxN_0__in_data_50),
    .in_data_51(muxN_0__in_data_51),
    .in_data_52(muxN_0__in_data_52),
    .in_data_53(muxN_0__in_data_53),
    .in_data_54(muxN_0__in_data_54),
    .in_data_55(muxN_0__in_data_55),
    .in_data_56(muxN_0__in_data_56),
    .in_data_57(muxN_0__in_data_57),
    .in_data_58(muxN_0__in_data_58),
    .in_data_59(muxN_0__in_data_59),
    .in_data_6(muxN_0__in_data_6),
    .in_data_60(muxN_0__in_data_60),
    .in_data_61(muxN_0__in_data_61),
    .in_data_62(muxN_0__in_data_62),
    .in_data_63(muxN_0__in_data_63),
    .in_data_7(muxN_0__in_data_7),
    .in_data_8(muxN_0__in_data_8),
    .in_data_9(muxN_0__in_data_9),
    .in_sel(muxN_0__in_sel),
    .out(muxN_0__out)
  );

  // Instancing generated Module: commonlib.muxn(N:16, width:32)
  wire [31:0] muxN_1__in_data_0;
  wire [31:0] muxN_1__in_data_1;
  wire [31:0] muxN_1__in_data_10;
  wire [31:0] muxN_1__in_data_11;
  wire [31:0] muxN_1__in_data_12;
  wire [31:0] muxN_1__in_data_13;
  wire [31:0] muxN_1__in_data_14;
  wire [31:0] muxN_1__in_data_15;
  wire [31:0] muxN_1__in_data_2;
  wire [31:0] muxN_1__in_data_3;
  wire [31:0] muxN_1__in_data_4;
  wire [31:0] muxN_1__in_data_5;
  wire [31:0] muxN_1__in_data_6;
  wire [31:0] muxN_1__in_data_7;
  wire [31:0] muxN_1__in_data_8;
  wire [31:0] muxN_1__in_data_9;
  wire [3:0] muxN_1__in_sel;
  wire [31:0] muxN_1__out;
  commonlib_muxn__N16__width32 muxN_1(
    .in_data_0(muxN_1__in_data_0),
    .in_data_1(muxN_1__in_data_1),
    .in_data_10(muxN_1__in_data_10),
    .in_data_11(muxN_1__in_data_11),
    .in_data_12(muxN_1__in_data_12),
    .in_data_13(muxN_1__in_data_13),
    .in_data_14(muxN_1__in_data_14),
    .in_data_15(muxN_1__in_data_15),
    .in_data_2(muxN_1__in_data_2),
    .in_data_3(muxN_1__in_data_3),
    .in_data_4(muxN_1__in_data_4),
    .in_data_5(muxN_1__in_data_5),
    .in_data_6(muxN_1__in_data_6),
    .in_data_7(muxN_1__in_data_7),
    .in_data_8(muxN_1__in_data_8),
    .in_data_9(muxN_1__in_data_9),
    .in_sel(muxN_1__in_sel),
    .out(muxN_1__out)
  );

  // Instancing generated Module: coreir.slice(hi:6, lo:0, width:7)
  wire [6:0] sel_slice0__in;
  wire [5:0] sel_slice0__out;
  coreir_slice #(.hi(6),.lo(0),.width(7)) sel_slice0(
    .in(sel_slice0__in),
    .out(sel_slice0__out)
  );

  // Instancing generated Module: coreir.slice(hi:4, lo:0, width:7)
  wire [6:0] sel_slice1__in;
  wire [3:0] sel_slice1__out;
  coreir_slice #(.hi(4),.lo(0),.width(7)) sel_slice1(
    .in(sel_slice1__in),
    .out(sel_slice1__out)
  );

  assign _join__in0[31:0] = muxN_0__out[31:0];

  assign _join__in1[31:0] = muxN_1__out[31:0];

  assign out[31:0] = _join__out[31:0];

  assign _join__sel = in_sel[6];

  assign muxN_0__in_data_0[31:0] = in_data_0[31:0];

  assign muxN_0__in_data_1[31:0] = in_data_1[31:0];

  assign muxN_0__in_data_10[31:0] = in_data_10[31:0];

  assign muxN_0__in_data_11[31:0] = in_data_11[31:0];

  assign muxN_0__in_data_12[31:0] = in_data_12[31:0];

  assign muxN_0__in_data_13[31:0] = in_data_13[31:0];

  assign muxN_0__in_data_14[31:0] = in_data_14[31:0];

  assign muxN_0__in_data_15[31:0] = in_data_15[31:0];

  assign muxN_0__in_data_16[31:0] = in_data_16[31:0];

  assign muxN_0__in_data_17[31:0] = in_data_17[31:0];

  assign muxN_0__in_data_18[31:0] = in_data_18[31:0];

  assign muxN_0__in_data_19[31:0] = in_data_19[31:0];

  assign muxN_0__in_data_2[31:0] = in_data_2[31:0];

  assign muxN_0__in_data_20[31:0] = in_data_20[31:0];

  assign muxN_0__in_data_21[31:0] = in_data_21[31:0];

  assign muxN_0__in_data_22[31:0] = in_data_22[31:0];

  assign muxN_0__in_data_23[31:0] = in_data_23[31:0];

  assign muxN_0__in_data_24[31:0] = in_data_24[31:0];

  assign muxN_0__in_data_25[31:0] = in_data_25[31:0];

  assign muxN_0__in_data_26[31:0] = in_data_26[31:0];

  assign muxN_0__in_data_27[31:0] = in_data_27[31:0];

  assign muxN_0__in_data_28[31:0] = in_data_28[31:0];

  assign muxN_0__in_data_29[31:0] = in_data_29[31:0];

  assign muxN_0__in_data_3[31:0] = in_data_3[31:0];

  assign muxN_0__in_data_30[31:0] = in_data_30[31:0];

  assign muxN_0__in_data_31[31:0] = in_data_31[31:0];

  assign muxN_0__in_data_32[31:0] = in_data_32[31:0];

  assign muxN_0__in_data_33[31:0] = in_data_33[31:0];

  assign muxN_0__in_data_34[31:0] = in_data_34[31:0];

  assign muxN_0__in_data_35[31:0] = in_data_35[31:0];

  assign muxN_0__in_data_36[31:0] = in_data_36[31:0];

  assign muxN_0__in_data_37[31:0] = in_data_37[31:0];

  assign muxN_0__in_data_38[31:0] = in_data_38[31:0];

  assign muxN_0__in_data_39[31:0] = in_data_39[31:0];

  assign muxN_0__in_data_4[31:0] = in_data_4[31:0];

  assign muxN_0__in_data_40[31:0] = in_data_40[31:0];

  assign muxN_0__in_data_41[31:0] = in_data_41[31:0];

  assign muxN_0__in_data_42[31:0] = in_data_42[31:0];

  assign muxN_0__in_data_43[31:0] = in_data_43[31:0];

  assign muxN_0__in_data_44[31:0] = in_data_44[31:0];

  assign muxN_0__in_data_45[31:0] = in_data_45[31:0];

  assign muxN_0__in_data_46[31:0] = in_data_46[31:0];

  assign muxN_0__in_data_47[31:0] = in_data_47[31:0];

  assign muxN_0__in_data_48[31:0] = in_data_48[31:0];

  assign muxN_0__in_data_49[31:0] = in_data_49[31:0];

  assign muxN_0__in_data_5[31:0] = in_data_5[31:0];

  assign muxN_0__in_data_50[31:0] = in_data_50[31:0];

  assign muxN_0__in_data_51[31:0] = in_data_51[31:0];

  assign muxN_0__in_data_52[31:0] = in_data_52[31:0];

  assign muxN_0__in_data_53[31:0] = in_data_53[31:0];

  assign muxN_0__in_data_54[31:0] = in_data_54[31:0];

  assign muxN_0__in_data_55[31:0] = in_data_55[31:0];

  assign muxN_0__in_data_56[31:0] = in_data_56[31:0];

  assign muxN_0__in_data_57[31:0] = in_data_57[31:0];

  assign muxN_0__in_data_58[31:0] = in_data_58[31:0];

  assign muxN_0__in_data_59[31:0] = in_data_59[31:0];

  assign muxN_0__in_data_6[31:0] = in_data_6[31:0];

  assign muxN_0__in_data_60[31:0] = in_data_60[31:0];

  assign muxN_0__in_data_61[31:0] = in_data_61[31:0];

  assign muxN_0__in_data_62[31:0] = in_data_62[31:0];

  assign muxN_0__in_data_63[31:0] = in_data_63[31:0];

  assign muxN_0__in_data_7[31:0] = in_data_7[31:0];

  assign muxN_0__in_data_8[31:0] = in_data_8[31:0];

  assign muxN_0__in_data_9[31:0] = in_data_9[31:0];

  assign muxN_0__in_sel[5:0] = sel_slice0__out[5:0];

  assign muxN_1__in_data_0[31:0] = in_data_64[31:0];

  assign muxN_1__in_data_1[31:0] = in_data_65[31:0];

  assign muxN_1__in_data_10[31:0] = in_data_74[31:0];

  assign muxN_1__in_data_11[31:0] = in_data_75[31:0];

  assign muxN_1__in_data_12[31:0] = in_data_76[31:0];

  assign muxN_1__in_data_13[31:0] = in_data_77[31:0];

  assign muxN_1__in_data_14[31:0] = in_data_78[31:0];

  assign muxN_1__in_data_15[31:0] = in_data_79[31:0];

  assign muxN_1__in_data_2[31:0] = in_data_66[31:0];

  assign muxN_1__in_data_3[31:0] = in_data_67[31:0];

  assign muxN_1__in_data_4[31:0] = in_data_68[31:0];

  assign muxN_1__in_data_5[31:0] = in_data_69[31:0];

  assign muxN_1__in_data_6[31:0] = in_data_70[31:0];

  assign muxN_1__in_data_7[31:0] = in_data_71[31:0];

  assign muxN_1__in_data_8[31:0] = in_data_72[31:0];

  assign muxN_1__in_data_9[31:0] = in_data_73[31:0];

  assign muxN_1__in_sel[3:0] = sel_slice1__out[3:0];

  assign sel_slice0__in[6:0] = in_sel[6:0];

  assign sel_slice1__in[6:0] = in_sel[6:0];


endmodule  // commonlib_muxn__N80__width32

// Generated from commonlib.muxn(N:10, width:16)
module commonlib_muxn__N10__width16 (
  input [15:0] in_data_0,
  input [15:0] in_data_1,
  input [15:0] in_data_2,
  input [15:0] in_data_3,
  input [15:0] in_data_4,
  input [15:0] in_data_5,
  input [15:0] in_data_6,
  input [15:0] in_data_7,
  input [15:0] in_data_8,
  input [15:0] in_data_9,
  input [3:0] in_sel,
  output [15:0] out
);


  // Instancing generated Module: coreir.mux(width:16)
  wire [15:0] _join__in0;
  wire [15:0] _join__in1;
  wire [15:0] _join__out;
  wire  _join__sel;
  coreir_mux #(.width(16)) _join(
    .in0(_join__in0),
    .in1(_join__in1),
    .out(_join__out),
    .sel(_join__sel)
  );

  // Instancing generated Module: commonlib.muxn(N:8, width:16)
  wire [15:0] muxN_0__in_data_0;
  wire [15:0] muxN_0__in_data_1;
  wire [15:0] muxN_0__in_data_2;
  wire [15:0] muxN_0__in_data_3;
  wire [15:0] muxN_0__in_data_4;
  wire [15:0] muxN_0__in_data_5;
  wire [15:0] muxN_0__in_data_6;
  wire [15:0] muxN_0__in_data_7;
  wire [2:0] muxN_0__in_sel;
  wire [15:0] muxN_0__out;
  commonlib_muxn__N8__width16 muxN_0(
    .in_data_0(muxN_0__in_data_0),
    .in_data_1(muxN_0__in_data_1),
    .in_data_2(muxN_0__in_data_2),
    .in_data_3(muxN_0__in_data_3),
    .in_data_4(muxN_0__in_data_4),
    .in_data_5(muxN_0__in_data_5),
    .in_data_6(muxN_0__in_data_6),
    .in_data_7(muxN_0__in_data_7),
    .in_sel(muxN_0__in_sel),
    .out(muxN_0__out)
  );

  // Instancing generated Module: commonlib.muxn(N:2, width:16)
  wire [15:0] muxN_1__in_data_0;
  wire [15:0] muxN_1__in_data_1;
  wire [0:0] muxN_1__in_sel;
  wire [15:0] muxN_1__out;
  commonlib_muxn__N2__width16 muxN_1(
    .in_data_0(muxN_1__in_data_0),
    .in_data_1(muxN_1__in_data_1),
    .in_sel(muxN_1__in_sel),
    .out(muxN_1__out)
  );

  // Instancing generated Module: coreir.slice(hi:3, lo:0, width:4)
  wire [3:0] sel_slice0__in;
  wire [2:0] sel_slice0__out;
  coreir_slice #(.hi(3),.lo(0),.width(4)) sel_slice0(
    .in(sel_slice0__in),
    .out(sel_slice0__out)
  );

  // Instancing generated Module: coreir.slice(hi:1, lo:0, width:4)
  wire [3:0] sel_slice1__in;
  wire [0:0] sel_slice1__out;
  coreir_slice #(.hi(1),.lo(0),.width(4)) sel_slice1(
    .in(sel_slice1__in),
    .out(sel_slice1__out)
  );

  assign _join__in0[15:0] = muxN_0__out[15:0];

  assign _join__in1[15:0] = muxN_1__out[15:0];

  assign out[15:0] = _join__out[15:0];

  assign _join__sel = in_sel[3];

  assign muxN_0__in_data_0[15:0] = in_data_0[15:0];

  assign muxN_0__in_data_1[15:0] = in_data_1[15:0];

  assign muxN_0__in_data_2[15:0] = in_data_2[15:0];

  assign muxN_0__in_data_3[15:0] = in_data_3[15:0];

  assign muxN_0__in_data_4[15:0] = in_data_4[15:0];

  assign muxN_0__in_data_5[15:0] = in_data_5[15:0];

  assign muxN_0__in_data_6[15:0] = in_data_6[15:0];

  assign muxN_0__in_data_7[15:0] = in_data_7[15:0];

  assign muxN_0__in_sel[2:0] = sel_slice0__out[2:0];

  assign muxN_1__in_data_0[15:0] = in_data_8[15:0];

  assign muxN_1__in_data_1[15:0] = in_data_9[15:0];

  assign muxN_1__in_sel[0:0] = sel_slice1__out[0:0];

  assign sel_slice0__in[3:0] = in_sel[3:0];

  assign sel_slice1__in[3:0] = in_sel[3:0];


endmodule  // commonlib_muxn__N10__width16

// Generated from commonlib.muxn(N:10, width:1)
module commonlib_muxn__N10__width1 (
  input [0:0] in_data_0,
  input [0:0] in_data_1,
  input [0:0] in_data_2,
  input [0:0] in_data_3,
  input [0:0] in_data_4,
  input [0:0] in_data_5,
  input [0:0] in_data_6,
  input [0:0] in_data_7,
  input [0:0] in_data_8,
  input [0:0] in_data_9,
  input [3:0] in_sel,
  output [0:0] out
);


  // Instancing generated Module: coreir.mux(width:1)
  wire [0:0] _join__in0;
  wire [0:0] _join__in1;
  wire [0:0] _join__out;
  wire  _join__sel;
  coreir_mux #(.width(1)) _join(
    .in0(_join__in0),
    .in1(_join__in1),
    .out(_join__out),
    .sel(_join__sel)
  );

  // Instancing generated Module: commonlib.muxn(N:8, width:1)
  wire [0:0] muxN_0__in_data_0;
  wire [0:0] muxN_0__in_data_1;
  wire [0:0] muxN_0__in_data_2;
  wire [0:0] muxN_0__in_data_3;
  wire [0:0] muxN_0__in_data_4;
  wire [0:0] muxN_0__in_data_5;
  wire [0:0] muxN_0__in_data_6;
  wire [0:0] muxN_0__in_data_7;
  wire [2:0] muxN_0__in_sel;
  wire [0:0] muxN_0__out;
  commonlib_muxn__N8__width1 muxN_0(
    .in_data_0(muxN_0__in_data_0),
    .in_data_1(muxN_0__in_data_1),
    .in_data_2(muxN_0__in_data_2),
    .in_data_3(muxN_0__in_data_3),
    .in_data_4(muxN_0__in_data_4),
    .in_data_5(muxN_0__in_data_5),
    .in_data_6(muxN_0__in_data_6),
    .in_data_7(muxN_0__in_data_7),
    .in_sel(muxN_0__in_sel),
    .out(muxN_0__out)
  );

  // Instancing generated Module: commonlib.muxn(N:2, width:1)
  wire [0:0] muxN_1__in_data_0;
  wire [0:0] muxN_1__in_data_1;
  wire [0:0] muxN_1__in_sel;
  wire [0:0] muxN_1__out;
  commonlib_muxn__N2__width1 muxN_1(
    .in_data_0(muxN_1__in_data_0),
    .in_data_1(muxN_1__in_data_1),
    .in_sel(muxN_1__in_sel),
    .out(muxN_1__out)
  );

  // Instancing generated Module: coreir.slice(hi:3, lo:0, width:4)
  wire [3:0] sel_slice0__in;
  wire [2:0] sel_slice0__out;
  coreir_slice #(.hi(3),.lo(0),.width(4)) sel_slice0(
    .in(sel_slice0__in),
    .out(sel_slice0__out)
  );

  // Instancing generated Module: coreir.slice(hi:1, lo:0, width:4)
  wire [3:0] sel_slice1__in;
  wire [0:0] sel_slice1__out;
  coreir_slice #(.hi(1),.lo(0),.width(4)) sel_slice1(
    .in(sel_slice1__in),
    .out(sel_slice1__out)
  );

  assign _join__in0[0:0] = muxN_0__out[0:0];

  assign _join__in1[0:0] = muxN_1__out[0:0];

  assign out[0:0] = _join__out[0:0];

  assign _join__sel = in_sel[3];

  assign muxN_0__in_data_0[0:0] = in_data_0[0:0];

  assign muxN_0__in_data_1[0:0] = in_data_1[0:0];

  assign muxN_0__in_data_2[0:0] = in_data_2[0:0];

  assign muxN_0__in_data_3[0:0] = in_data_3[0:0];

  assign muxN_0__in_data_4[0:0] = in_data_4[0:0];

  assign muxN_0__in_data_5[0:0] = in_data_5[0:0];

  assign muxN_0__in_data_6[0:0] = in_data_6[0:0];

  assign muxN_0__in_data_7[0:0] = in_data_7[0:0];

  assign muxN_0__in_sel[2:0] = sel_slice0__out[2:0];

  assign muxN_1__in_data_0[0:0] = in_data_8[0:0];

  assign muxN_1__in_data_1[0:0] = in_data_9[0:0];

  assign muxN_1__in_sel[0:0] = sel_slice1__out[0:0];

  assign sel_slice0__in[3:0] = in_sel[3:0];

  assign sel_slice1__in[3:0] = in_sel[3:0];


endmodule  // commonlib_muxn__N10__width1

module ZextWrapper_4_32 (
  input [3:0] I,
  output [31:0] O
);


  wire  bit_const_0_None__out;
  corebit_const #(.value(0)) bit_const_0_None(
    .out(bit_const_0_None__out)
  );

  assign O[10] = bit_const_0_None__out;

  assign O[11] = bit_const_0_None__out;

  assign O[12] = bit_const_0_None__out;

  assign O[13] = bit_const_0_None__out;

  assign O[14] = bit_const_0_None__out;

  assign O[15] = bit_const_0_None__out;

  assign O[16] = bit_const_0_None__out;

  assign O[17] = bit_const_0_None__out;

  assign O[18] = bit_const_0_None__out;

  assign O[19] = bit_const_0_None__out;

  assign O[20] = bit_const_0_None__out;

  assign O[21] = bit_const_0_None__out;

  assign O[22] = bit_const_0_None__out;

  assign O[23] = bit_const_0_None__out;

  assign O[24] = bit_const_0_None__out;

  assign O[25] = bit_const_0_None__out;

  assign O[26] = bit_const_0_None__out;

  assign O[27] = bit_const_0_None__out;

  assign O[28] = bit_const_0_None__out;

  assign O[29] = bit_const_0_None__out;

  assign O[30] = bit_const_0_None__out;

  assign O[31] = bit_const_0_None__out;

  assign O[4] = bit_const_0_None__out;

  assign O[5] = bit_const_0_None__out;

  assign O[6] = bit_const_0_None__out;

  assign O[7] = bit_const_0_None__out;

  assign O[8] = bit_const_0_None__out;

  assign O[9] = bit_const_0_None__out;

  assign O[0] = I[0];

  assign O[1] = I[1];

  assign O[2] = I[2];

  assign O[3] = I[3];


endmodule  // ZextWrapper_4_32

module ZextWrapper_2_32 (
  input [1:0] I,
  output [31:0] O
);


  wire  bit_const_0_None__out;
  corebit_const #(.value(0)) bit_const_0_None(
    .out(bit_const_0_None__out)
  );

  assign O[10] = bit_const_0_None__out;

  assign O[11] = bit_const_0_None__out;

  assign O[12] = bit_const_0_None__out;

  assign O[13] = bit_const_0_None__out;

  assign O[14] = bit_const_0_None__out;

  assign O[15] = bit_const_0_None__out;

  assign O[16] = bit_const_0_None__out;

  assign O[17] = bit_const_0_None__out;

  assign O[18] = bit_const_0_None__out;

  assign O[19] = bit_const_0_None__out;

  assign O[20] = bit_const_0_None__out;

  assign O[21] = bit_const_0_None__out;

  assign O[22] = bit_const_0_None__out;

  assign O[23] = bit_const_0_None__out;

  assign O[24] = bit_const_0_None__out;

  assign O[25] = bit_const_0_None__out;

  assign O[26] = bit_const_0_None__out;

  assign O[27] = bit_const_0_None__out;

  assign O[28] = bit_const_0_None__out;

  assign O[29] = bit_const_0_None__out;

  assign O[2] = bit_const_0_None__out;

  assign O[30] = bit_const_0_None__out;

  assign O[31] = bit_const_0_None__out;

  assign O[3] = bit_const_0_None__out;

  assign O[4] = bit_const_0_None__out;

  assign O[5] = bit_const_0_None__out;

  assign O[6] = bit_const_0_None__out;

  assign O[7] = bit_const_0_None__out;

  assign O[8] = bit_const_0_None__out;

  assign O[9] = bit_const_0_None__out;

  assign O[0] = I[0];

  assign O[1] = I[1];


endmodule  // ZextWrapper_2_32

module ZextWrapper_1_32 (
  input [0:0] I,
  output [31:0] O
);


  wire  bit_const_0_None__out;
  corebit_const #(.value(0)) bit_const_0_None(
    .out(bit_const_0_None__out)
  );

  assign O[10] = bit_const_0_None__out;

  assign O[11] = bit_const_0_None__out;

  assign O[12] = bit_const_0_None__out;

  assign O[13] = bit_const_0_None__out;

  assign O[14] = bit_const_0_None__out;

  assign O[15] = bit_const_0_None__out;

  assign O[16] = bit_const_0_None__out;

  assign O[17] = bit_const_0_None__out;

  assign O[18] = bit_const_0_None__out;

  assign O[19] = bit_const_0_None__out;

  assign O[1] = bit_const_0_None__out;

  assign O[20] = bit_const_0_None__out;

  assign O[21] = bit_const_0_None__out;

  assign O[22] = bit_const_0_None__out;

  assign O[23] = bit_const_0_None__out;

  assign O[24] = bit_const_0_None__out;

  assign O[25] = bit_const_0_None__out;

  assign O[26] = bit_const_0_None__out;

  assign O[27] = bit_const_0_None__out;

  assign O[28] = bit_const_0_None__out;

  assign O[29] = bit_const_0_None__out;

  assign O[2] = bit_const_0_None__out;

  assign O[30] = bit_const_0_None__out;

  assign O[31] = bit_const_0_None__out;

  assign O[3] = bit_const_0_None__out;

  assign O[4] = bit_const_0_None__out;

  assign O[5] = bit_const_0_None__out;

  assign O[6] = bit_const_0_None__out;

  assign O[7] = bit_const_0_None__out;

  assign O[8] = bit_const_0_None__out;

  assign O[9] = bit_const_0_None__out;

  assign O[0] = I[0];


endmodule  // ZextWrapper_1_32

module PECore (
  input [0:0] bit0,
  input [0:0] bit1,
  input [0:0] bit2,
  input  clk,
  input [7:0] config_config_addr,
  input [31:0] config_config_data,
  input [0:0] config_read,
  input [0:0] config_write,
  input [15:0] data0,
  input [15:0] data1,
  output [31:0] read_config_data,
  output [15:0] res,
  output [0:0] res_p,
  input  reset,
  input [3:0] stall
);


  // Instancing generated Module: coreir.not(width:1)
  wire [0:0] Invert1_inst0__in;
  wire [0:0] Invert1_inst0__out;
  coreir_not #(.width(1)) Invert1_inst0(
    .in(Invert1_inst0__in),
    .out(Invert1_inst0__out)
  );

  wire  test_pe_inst0__bit0;
  wire  test_pe_inst0__bit1;
  wire  test_pe_inst0__bit2;
  wire [7:0] test_pe_inst0__cfg_a;
  wire [31:0] test_pe_inst0__cfg_d;
  wire  test_pe_inst0__cfg_en;
  wire  test_pe_inst0__clk;
  wire  test_pe_inst0__clk_en;
  wire [15:0] test_pe_inst0__data0;
  wire [15:0] test_pe_inst0__data1;
  wire  test_pe_inst0__irq;
  wire [31:0] test_pe_inst0__read_data;
  wire [15:0] test_pe_inst0__res;
  wire  test_pe_inst0__res_p;
  wire  test_pe_inst0__rst_n;
  test_pe test_pe_inst0(
    .bit0(test_pe_inst0__bit0),
    .bit1(test_pe_inst0__bit1),
    .bit2(test_pe_inst0__bit2),
    .cfg_a(test_pe_inst0__cfg_a),
    .cfg_d(test_pe_inst0__cfg_d),
    .cfg_en(test_pe_inst0__cfg_en),
    .clk(test_pe_inst0__clk),
    .clk_en(test_pe_inst0__clk_en),
    .data0(test_pe_inst0__data0),
    .data1(test_pe_inst0__data1),
    .irq(test_pe_inst0__irq),
    .read_data(test_pe_inst0__read_data),
    .res(test_pe_inst0__res),
    .res_p(test_pe_inst0__res_p),
    .rst_n(test_pe_inst0__rst_n)
  );

  assign Invert1_inst0__in[0] = stall[0];

  assign test_pe_inst0__clk_en = Invert1_inst0__out[0];

  assign test_pe_inst0__bit0 = bit0[0];

  assign test_pe_inst0__bit1 = bit1[0];

  assign test_pe_inst0__bit2 = bit2[0];

  assign test_pe_inst0__clk = clk;

  assign test_pe_inst0__cfg_a[7:0] = config_config_addr[7:0];

  assign test_pe_inst0__cfg_d[31:0] = config_config_data[31:0];

  assign test_pe_inst0__cfg_en = config_write[0];

  assign test_pe_inst0__data0[15:0] = data0[15:0];

  assign test_pe_inst0__data1[15:0] = data1[15:0];

  assign read_config_data[31:0] = test_pe_inst0__read_data[31:0];

  assign res[15:0] = test_pe_inst0__res[15:0];

  assign res_p[0] = test_pe_inst0__res_p;

  assign test_pe_inst0__rst_n = reset;


endmodule  // PECore

module Mux80x32 (
  input [31:0] I0,
  input [31:0] I1,
  input [31:0] I10,
  input [31:0] I11,
  input [31:0] I12,
  input [31:0] I13,
  input [31:0] I14,
  input [31:0] I15,
  input [31:0] I16,
  input [31:0] I17,
  input [31:0] I18,
  input [31:0] I19,
  input [31:0] I2,
  input [31:0] I20,
  input [31:0] I21,
  input [31:0] I22,
  input [31:0] I23,
  input [31:0] I24,
  input [31:0] I25,
  input [31:0] I26,
  input [31:0] I27,
  input [31:0] I28,
  input [31:0] I29,
  input [31:0] I3,
  input [31:0] I30,
  input [31:0] I31,
  input [31:0] I32,
  input [31:0] I33,
  input [31:0] I34,
  input [31:0] I35,
  input [31:0] I36,
  input [31:0] I37,
  input [31:0] I38,
  input [31:0] I39,
  input [31:0] I4,
  input [31:0] I40,
  input [31:0] I41,
  input [31:0] I42,
  input [31:0] I43,
  input [31:0] I44,
  input [31:0] I45,
  input [31:0] I46,
  input [31:0] I47,
  input [31:0] I48,
  input [31:0] I49,
  input [31:0] I5,
  input [31:0] I50,
  input [31:0] I51,
  input [31:0] I52,
  input [31:0] I53,
  input [31:0] I54,
  input [31:0] I55,
  input [31:0] I56,
  input [31:0] I57,
  input [31:0] I58,
  input [31:0] I59,
  input [31:0] I6,
  input [31:0] I60,
  input [31:0] I61,
  input [31:0] I62,
  input [31:0] I63,
  input [31:0] I64,
  input [31:0] I65,
  input [31:0] I66,
  input [31:0] I67,
  input [31:0] I68,
  input [31:0] I69,
  input [31:0] I7,
  input [31:0] I70,
  input [31:0] I71,
  input [31:0] I72,
  input [31:0] I73,
  input [31:0] I74,
  input [31:0] I75,
  input [31:0] I76,
  input [31:0] I77,
  input [31:0] I78,
  input [31:0] I79,
  input [31:0] I8,
  input [31:0] I9,
  output [31:0] O,
  input [6:0] S
);


  // Instancing generated Module: commonlib.muxn(N:80, width:32)
  wire [31:0] coreir_commonlib_mux80x32_inst0__in_data_0;
  wire [31:0] coreir_commonlib_mux80x32_inst0__in_data_1;
  wire [31:0] coreir_commonlib_mux80x32_inst0__in_data_10;
  wire [31:0] coreir_commonlib_mux80x32_inst0__in_data_11;
  wire [31:0] coreir_commonlib_mux80x32_inst0__in_data_12;
  wire [31:0] coreir_commonlib_mux80x32_inst0__in_data_13;
  wire [31:0] coreir_commonlib_mux80x32_inst0__in_data_14;
  wire [31:0] coreir_commonlib_mux80x32_inst0__in_data_15;
  wire [31:0] coreir_commonlib_mux80x32_inst0__in_data_16;
  wire [31:0] coreir_commonlib_mux80x32_inst0__in_data_17;
  wire [31:0] coreir_commonlib_mux80x32_inst0__in_data_18;
  wire [31:0] coreir_commonlib_mux80x32_inst0__in_data_19;
  wire [31:0] coreir_commonlib_mux80x32_inst0__in_data_2;
  wire [31:0] coreir_commonlib_mux80x32_inst0__in_data_20;
  wire [31:0] coreir_commonlib_mux80x32_inst0__in_data_21;
  wire [31:0] coreir_commonlib_mux80x32_inst0__in_data_22;
  wire [31:0] coreir_commonlib_mux80x32_inst0__in_data_23;
  wire [31:0] coreir_commonlib_mux80x32_inst0__in_data_24;
  wire [31:0] coreir_commonlib_mux80x32_inst0__in_data_25;
  wire [31:0] coreir_commonlib_mux80x32_inst0__in_data_26;
  wire [31:0] coreir_commonlib_mux80x32_inst0__in_data_27;
  wire [31:0] coreir_commonlib_mux80x32_inst0__in_data_28;
  wire [31:0] coreir_commonlib_mux80x32_inst0__in_data_29;
  wire [31:0] coreir_commonlib_mux80x32_inst0__in_data_3;
  wire [31:0] coreir_commonlib_mux80x32_inst0__in_data_30;
  wire [31:0] coreir_commonlib_mux80x32_inst0__in_data_31;
  wire [31:0] coreir_commonlib_mux80x32_inst0__in_data_32;
  wire [31:0] coreir_commonlib_mux80x32_inst0__in_data_33;
  wire [31:0] coreir_commonlib_mux80x32_inst0__in_data_34;
  wire [31:0] coreir_commonlib_mux80x32_inst0__in_data_35;
  wire [31:0] coreir_commonlib_mux80x32_inst0__in_data_36;
  wire [31:0] coreir_commonlib_mux80x32_inst0__in_data_37;
  wire [31:0] coreir_commonlib_mux80x32_inst0__in_data_38;
  wire [31:0] coreir_commonlib_mux80x32_inst0__in_data_39;
  wire [31:0] coreir_commonlib_mux80x32_inst0__in_data_4;
  wire [31:0] coreir_commonlib_mux80x32_inst0__in_data_40;
  wire [31:0] coreir_commonlib_mux80x32_inst0__in_data_41;
  wire [31:0] coreir_commonlib_mux80x32_inst0__in_data_42;
  wire [31:0] coreir_commonlib_mux80x32_inst0__in_data_43;
  wire [31:0] coreir_commonlib_mux80x32_inst0__in_data_44;
  wire [31:0] coreir_commonlib_mux80x32_inst0__in_data_45;
  wire [31:0] coreir_commonlib_mux80x32_inst0__in_data_46;
  wire [31:0] coreir_commonlib_mux80x32_inst0__in_data_47;
  wire [31:0] coreir_commonlib_mux80x32_inst0__in_data_48;
  wire [31:0] coreir_commonlib_mux80x32_inst0__in_data_49;
  wire [31:0] coreir_commonlib_mux80x32_inst0__in_data_5;
  wire [31:0] coreir_commonlib_mux80x32_inst0__in_data_50;
  wire [31:0] coreir_commonlib_mux80x32_inst0__in_data_51;
  wire [31:0] coreir_commonlib_mux80x32_inst0__in_data_52;
  wire [31:0] coreir_commonlib_mux80x32_inst0__in_data_53;
  wire [31:0] coreir_commonlib_mux80x32_inst0__in_data_54;
  wire [31:0] coreir_commonlib_mux80x32_inst0__in_data_55;
  wire [31:0] coreir_commonlib_mux80x32_inst0__in_data_56;
  wire [31:0] coreir_commonlib_mux80x32_inst0__in_data_57;
  wire [31:0] coreir_commonlib_mux80x32_inst0__in_data_58;
  wire [31:0] coreir_commonlib_mux80x32_inst0__in_data_59;
  wire [31:0] coreir_commonlib_mux80x32_inst0__in_data_6;
  wire [31:0] coreir_commonlib_mux80x32_inst0__in_data_60;
  wire [31:0] coreir_commonlib_mux80x32_inst0__in_data_61;
  wire [31:0] coreir_commonlib_mux80x32_inst0__in_data_62;
  wire [31:0] coreir_commonlib_mux80x32_inst0__in_data_63;
  wire [31:0] coreir_commonlib_mux80x32_inst0__in_data_64;
  wire [31:0] coreir_commonlib_mux80x32_inst0__in_data_65;
  wire [31:0] coreir_commonlib_mux80x32_inst0__in_data_66;
  wire [31:0] coreir_commonlib_mux80x32_inst0__in_data_67;
  wire [31:0] coreir_commonlib_mux80x32_inst0__in_data_68;
  wire [31:0] coreir_commonlib_mux80x32_inst0__in_data_69;
  wire [31:0] coreir_commonlib_mux80x32_inst0__in_data_7;
  wire [31:0] coreir_commonlib_mux80x32_inst0__in_data_70;
  wire [31:0] coreir_commonlib_mux80x32_inst0__in_data_71;
  wire [31:0] coreir_commonlib_mux80x32_inst0__in_data_72;
  wire [31:0] coreir_commonlib_mux80x32_inst0__in_data_73;
  wire [31:0] coreir_commonlib_mux80x32_inst0__in_data_74;
  wire [31:0] coreir_commonlib_mux80x32_inst0__in_data_75;
  wire [31:0] coreir_commonlib_mux80x32_inst0__in_data_76;
  wire [31:0] coreir_commonlib_mux80x32_inst0__in_data_77;
  wire [31:0] coreir_commonlib_mux80x32_inst0__in_data_78;
  wire [31:0] coreir_commonlib_mux80x32_inst0__in_data_79;
  wire [31:0] coreir_commonlib_mux80x32_inst0__in_data_8;
  wire [31:0] coreir_commonlib_mux80x32_inst0__in_data_9;
  wire [6:0] coreir_commonlib_mux80x32_inst0__in_sel;
  wire [31:0] coreir_commonlib_mux80x32_inst0__out;
  commonlib_muxn__N80__width32 coreir_commonlib_mux80x32_inst0(
    .in_data_0(coreir_commonlib_mux80x32_inst0__in_data_0),
    .in_data_1(coreir_commonlib_mux80x32_inst0__in_data_1),
    .in_data_10(coreir_commonlib_mux80x32_inst0__in_data_10),
    .in_data_11(coreir_commonlib_mux80x32_inst0__in_data_11),
    .in_data_12(coreir_commonlib_mux80x32_inst0__in_data_12),
    .in_data_13(coreir_commonlib_mux80x32_inst0__in_data_13),
    .in_data_14(coreir_commonlib_mux80x32_inst0__in_data_14),
    .in_data_15(coreir_commonlib_mux80x32_inst0__in_data_15),
    .in_data_16(coreir_commonlib_mux80x32_inst0__in_data_16),
    .in_data_17(coreir_commonlib_mux80x32_inst0__in_data_17),
    .in_data_18(coreir_commonlib_mux80x32_inst0__in_data_18),
    .in_data_19(coreir_commonlib_mux80x32_inst0__in_data_19),
    .in_data_2(coreir_commonlib_mux80x32_inst0__in_data_2),
    .in_data_20(coreir_commonlib_mux80x32_inst0__in_data_20),
    .in_data_21(coreir_commonlib_mux80x32_inst0__in_data_21),
    .in_data_22(coreir_commonlib_mux80x32_inst0__in_data_22),
    .in_data_23(coreir_commonlib_mux80x32_inst0__in_data_23),
    .in_data_24(coreir_commonlib_mux80x32_inst0__in_data_24),
    .in_data_25(coreir_commonlib_mux80x32_inst0__in_data_25),
    .in_data_26(coreir_commonlib_mux80x32_inst0__in_data_26),
    .in_data_27(coreir_commonlib_mux80x32_inst0__in_data_27),
    .in_data_28(coreir_commonlib_mux80x32_inst0__in_data_28),
    .in_data_29(coreir_commonlib_mux80x32_inst0__in_data_29),
    .in_data_3(coreir_commonlib_mux80x32_inst0__in_data_3),
    .in_data_30(coreir_commonlib_mux80x32_inst0__in_data_30),
    .in_data_31(coreir_commonlib_mux80x32_inst0__in_data_31),
    .in_data_32(coreir_commonlib_mux80x32_inst0__in_data_32),
    .in_data_33(coreir_commonlib_mux80x32_inst0__in_data_33),
    .in_data_34(coreir_commonlib_mux80x32_inst0__in_data_34),
    .in_data_35(coreir_commonlib_mux80x32_inst0__in_data_35),
    .in_data_36(coreir_commonlib_mux80x32_inst0__in_data_36),
    .in_data_37(coreir_commonlib_mux80x32_inst0__in_data_37),
    .in_data_38(coreir_commonlib_mux80x32_inst0__in_data_38),
    .in_data_39(coreir_commonlib_mux80x32_inst0__in_data_39),
    .in_data_4(coreir_commonlib_mux80x32_inst0__in_data_4),
    .in_data_40(coreir_commonlib_mux80x32_inst0__in_data_40),
    .in_data_41(coreir_commonlib_mux80x32_inst0__in_data_41),
    .in_data_42(coreir_commonlib_mux80x32_inst0__in_data_42),
    .in_data_43(coreir_commonlib_mux80x32_inst0__in_data_43),
    .in_data_44(coreir_commonlib_mux80x32_inst0__in_data_44),
    .in_data_45(coreir_commonlib_mux80x32_inst0__in_data_45),
    .in_data_46(coreir_commonlib_mux80x32_inst0__in_data_46),
    .in_data_47(coreir_commonlib_mux80x32_inst0__in_data_47),
    .in_data_48(coreir_commonlib_mux80x32_inst0__in_data_48),
    .in_data_49(coreir_commonlib_mux80x32_inst0__in_data_49),
    .in_data_5(coreir_commonlib_mux80x32_inst0__in_data_5),
    .in_data_50(coreir_commonlib_mux80x32_inst0__in_data_50),
    .in_data_51(coreir_commonlib_mux80x32_inst0__in_data_51),
    .in_data_52(coreir_commonlib_mux80x32_inst0__in_data_52),
    .in_data_53(coreir_commonlib_mux80x32_inst0__in_data_53),
    .in_data_54(coreir_commonlib_mux80x32_inst0__in_data_54),
    .in_data_55(coreir_commonlib_mux80x32_inst0__in_data_55),
    .in_data_56(coreir_commonlib_mux80x32_inst0__in_data_56),
    .in_data_57(coreir_commonlib_mux80x32_inst0__in_data_57),
    .in_data_58(coreir_commonlib_mux80x32_inst0__in_data_58),
    .in_data_59(coreir_commonlib_mux80x32_inst0__in_data_59),
    .in_data_6(coreir_commonlib_mux80x32_inst0__in_data_6),
    .in_data_60(coreir_commonlib_mux80x32_inst0__in_data_60),
    .in_data_61(coreir_commonlib_mux80x32_inst0__in_data_61),
    .in_data_62(coreir_commonlib_mux80x32_inst0__in_data_62),
    .in_data_63(coreir_commonlib_mux80x32_inst0__in_data_63),
    .in_data_64(coreir_commonlib_mux80x32_inst0__in_data_64),
    .in_data_65(coreir_commonlib_mux80x32_inst0__in_data_65),
    .in_data_66(coreir_commonlib_mux80x32_inst0__in_data_66),
    .in_data_67(coreir_commonlib_mux80x32_inst0__in_data_67),
    .in_data_68(coreir_commonlib_mux80x32_inst0__in_data_68),
    .in_data_69(coreir_commonlib_mux80x32_inst0__in_data_69),
    .in_data_7(coreir_commonlib_mux80x32_inst0__in_data_7),
    .in_data_70(coreir_commonlib_mux80x32_inst0__in_data_70),
    .in_data_71(coreir_commonlib_mux80x32_inst0__in_data_71),
    .in_data_72(coreir_commonlib_mux80x32_inst0__in_data_72),
    .in_data_73(coreir_commonlib_mux80x32_inst0__in_data_73),
    .in_data_74(coreir_commonlib_mux80x32_inst0__in_data_74),
    .in_data_75(coreir_commonlib_mux80x32_inst0__in_data_75),
    .in_data_76(coreir_commonlib_mux80x32_inst0__in_data_76),
    .in_data_77(coreir_commonlib_mux80x32_inst0__in_data_77),
    .in_data_78(coreir_commonlib_mux80x32_inst0__in_data_78),
    .in_data_79(coreir_commonlib_mux80x32_inst0__in_data_79),
    .in_data_8(coreir_commonlib_mux80x32_inst0__in_data_8),
    .in_data_9(coreir_commonlib_mux80x32_inst0__in_data_9),
    .in_sel(coreir_commonlib_mux80x32_inst0__in_sel),
    .out(coreir_commonlib_mux80x32_inst0__out)
  );

  assign coreir_commonlib_mux80x32_inst0__in_data_0[31:0] = I0[31:0];

  assign coreir_commonlib_mux80x32_inst0__in_data_1[31:0] = I1[31:0];

  assign coreir_commonlib_mux80x32_inst0__in_data_10[31:0] = I10[31:0];

  assign coreir_commonlib_mux80x32_inst0__in_data_11[31:0] = I11[31:0];

  assign coreir_commonlib_mux80x32_inst0__in_data_12[31:0] = I12[31:0];

  assign coreir_commonlib_mux80x32_inst0__in_data_13[31:0] = I13[31:0];

  assign coreir_commonlib_mux80x32_inst0__in_data_14[31:0] = I14[31:0];

  assign coreir_commonlib_mux80x32_inst0__in_data_15[31:0] = I15[31:0];

  assign coreir_commonlib_mux80x32_inst0__in_data_16[31:0] = I16[31:0];

  assign coreir_commonlib_mux80x32_inst0__in_data_17[31:0] = I17[31:0];

  assign coreir_commonlib_mux80x32_inst0__in_data_18[31:0] = I18[31:0];

  assign coreir_commonlib_mux80x32_inst0__in_data_19[31:0] = I19[31:0];

  assign coreir_commonlib_mux80x32_inst0__in_data_2[31:0] = I2[31:0];

  assign coreir_commonlib_mux80x32_inst0__in_data_20[31:0] = I20[31:0];

  assign coreir_commonlib_mux80x32_inst0__in_data_21[31:0] = I21[31:0];

  assign coreir_commonlib_mux80x32_inst0__in_data_22[31:0] = I22[31:0];

  assign coreir_commonlib_mux80x32_inst0__in_data_23[31:0] = I23[31:0];

  assign coreir_commonlib_mux80x32_inst0__in_data_24[31:0] = I24[31:0];

  assign coreir_commonlib_mux80x32_inst0__in_data_25[31:0] = I25[31:0];

  assign coreir_commonlib_mux80x32_inst0__in_data_26[31:0] = I26[31:0];

  assign coreir_commonlib_mux80x32_inst0__in_data_27[31:0] = I27[31:0];

  assign coreir_commonlib_mux80x32_inst0__in_data_28[31:0] = I28[31:0];

  assign coreir_commonlib_mux80x32_inst0__in_data_29[31:0] = I29[31:0];

  assign coreir_commonlib_mux80x32_inst0__in_data_3[31:0] = I3[31:0];

  assign coreir_commonlib_mux80x32_inst0__in_data_30[31:0] = I30[31:0];

  assign coreir_commonlib_mux80x32_inst0__in_data_31[31:0] = I31[31:0];

  assign coreir_commonlib_mux80x32_inst0__in_data_32[31:0] = I32[31:0];

  assign coreir_commonlib_mux80x32_inst0__in_data_33[31:0] = I33[31:0];

  assign coreir_commonlib_mux80x32_inst0__in_data_34[31:0] = I34[31:0];

  assign coreir_commonlib_mux80x32_inst0__in_data_35[31:0] = I35[31:0];

  assign coreir_commonlib_mux80x32_inst0__in_data_36[31:0] = I36[31:0];

  assign coreir_commonlib_mux80x32_inst0__in_data_37[31:0] = I37[31:0];

  assign coreir_commonlib_mux80x32_inst0__in_data_38[31:0] = I38[31:0];

  assign coreir_commonlib_mux80x32_inst0__in_data_39[31:0] = I39[31:0];

  assign coreir_commonlib_mux80x32_inst0__in_data_4[31:0] = I4[31:0];

  assign coreir_commonlib_mux80x32_inst0__in_data_40[31:0] = I40[31:0];

  assign coreir_commonlib_mux80x32_inst0__in_data_41[31:0] = I41[31:0];

  assign coreir_commonlib_mux80x32_inst0__in_data_42[31:0] = I42[31:0];

  assign coreir_commonlib_mux80x32_inst0__in_data_43[31:0] = I43[31:0];

  assign coreir_commonlib_mux80x32_inst0__in_data_44[31:0] = I44[31:0];

  assign coreir_commonlib_mux80x32_inst0__in_data_45[31:0] = I45[31:0];

  assign coreir_commonlib_mux80x32_inst0__in_data_46[31:0] = I46[31:0];

  assign coreir_commonlib_mux80x32_inst0__in_data_47[31:0] = I47[31:0];

  assign coreir_commonlib_mux80x32_inst0__in_data_48[31:0] = I48[31:0];

  assign coreir_commonlib_mux80x32_inst0__in_data_49[31:0] = I49[31:0];

  assign coreir_commonlib_mux80x32_inst0__in_data_5[31:0] = I5[31:0];

  assign coreir_commonlib_mux80x32_inst0__in_data_50[31:0] = I50[31:0];

  assign coreir_commonlib_mux80x32_inst0__in_data_51[31:0] = I51[31:0];

  assign coreir_commonlib_mux80x32_inst0__in_data_52[31:0] = I52[31:0];

  assign coreir_commonlib_mux80x32_inst0__in_data_53[31:0] = I53[31:0];

  assign coreir_commonlib_mux80x32_inst0__in_data_54[31:0] = I54[31:0];

  assign coreir_commonlib_mux80x32_inst0__in_data_55[31:0] = I55[31:0];

  assign coreir_commonlib_mux80x32_inst0__in_data_56[31:0] = I56[31:0];

  assign coreir_commonlib_mux80x32_inst0__in_data_57[31:0] = I57[31:0];

  assign coreir_commonlib_mux80x32_inst0__in_data_58[31:0] = I58[31:0];

  assign coreir_commonlib_mux80x32_inst0__in_data_59[31:0] = I59[31:0];

  assign coreir_commonlib_mux80x32_inst0__in_data_6[31:0] = I6[31:0];

  assign coreir_commonlib_mux80x32_inst0__in_data_60[31:0] = I60[31:0];

  assign coreir_commonlib_mux80x32_inst0__in_data_61[31:0] = I61[31:0];

  assign coreir_commonlib_mux80x32_inst0__in_data_62[31:0] = I62[31:0];

  assign coreir_commonlib_mux80x32_inst0__in_data_63[31:0] = I63[31:0];

  assign coreir_commonlib_mux80x32_inst0__in_data_64[31:0] = I64[31:0];

  assign coreir_commonlib_mux80x32_inst0__in_data_65[31:0] = I65[31:0];

  assign coreir_commonlib_mux80x32_inst0__in_data_66[31:0] = I66[31:0];

  assign coreir_commonlib_mux80x32_inst0__in_data_67[31:0] = I67[31:0];

  assign coreir_commonlib_mux80x32_inst0__in_data_68[31:0] = I68[31:0];

  assign coreir_commonlib_mux80x32_inst0__in_data_69[31:0] = I69[31:0];

  assign coreir_commonlib_mux80x32_inst0__in_data_7[31:0] = I7[31:0];

  assign coreir_commonlib_mux80x32_inst0__in_data_70[31:0] = I70[31:0];

  assign coreir_commonlib_mux80x32_inst0__in_data_71[31:0] = I71[31:0];

  assign coreir_commonlib_mux80x32_inst0__in_data_72[31:0] = I72[31:0];

  assign coreir_commonlib_mux80x32_inst0__in_data_73[31:0] = I73[31:0];

  assign coreir_commonlib_mux80x32_inst0__in_data_74[31:0] = I74[31:0];

  assign coreir_commonlib_mux80x32_inst0__in_data_75[31:0] = I75[31:0];

  assign coreir_commonlib_mux80x32_inst0__in_data_76[31:0] = I76[31:0];

  assign coreir_commonlib_mux80x32_inst0__in_data_77[31:0] = I77[31:0];

  assign coreir_commonlib_mux80x32_inst0__in_data_78[31:0] = I78[31:0];

  assign coreir_commonlib_mux80x32_inst0__in_data_79[31:0] = I79[31:0];

  assign coreir_commonlib_mux80x32_inst0__in_data_8[31:0] = I8[31:0];

  assign coreir_commonlib_mux80x32_inst0__in_data_9[31:0] = I9[31:0];

  assign coreir_commonlib_mux80x32_inst0__in_sel[6:0] = S[6:0];

  assign O[31:0] = coreir_commonlib_mux80x32_inst0__out[31:0];


endmodule  // Mux80x32

module MuxWrapper_80_32 (
  input [31:0] I_0,
  input [31:0] I_1,
  input [31:0] I_10,
  input [31:0] I_11,
  input [31:0] I_12,
  input [31:0] I_13,
  input [31:0] I_14,
  input [31:0] I_15,
  input [31:0] I_16,
  input [31:0] I_17,
  input [31:0] I_18,
  input [31:0] I_19,
  input [31:0] I_2,
  input [31:0] I_20,
  input [31:0] I_21,
  input [31:0] I_22,
  input [31:0] I_23,
  input [31:0] I_24,
  input [31:0] I_25,
  input [31:0] I_26,
  input [31:0] I_27,
  input [31:0] I_28,
  input [31:0] I_29,
  input [31:0] I_3,
  input [31:0] I_30,
  input [31:0] I_31,
  input [31:0] I_32,
  input [31:0] I_33,
  input [31:0] I_34,
  input [31:0] I_35,
  input [31:0] I_36,
  input [31:0] I_37,
  input [31:0] I_38,
  input [31:0] I_39,
  input [31:0] I_4,
  input [31:0] I_40,
  input [31:0] I_41,
  input [31:0] I_42,
  input [31:0] I_43,
  input [31:0] I_44,
  input [31:0] I_45,
  input [31:0] I_46,
  input [31:0] I_47,
  input [31:0] I_48,
  input [31:0] I_49,
  input [31:0] I_5,
  input [31:0] I_50,
  input [31:0] I_51,
  input [31:0] I_52,
  input [31:0] I_53,
  input [31:0] I_54,
  input [31:0] I_55,
  input [31:0] I_56,
  input [31:0] I_57,
  input [31:0] I_58,
  input [31:0] I_59,
  input [31:0] I_6,
  input [31:0] I_60,
  input [31:0] I_61,
  input [31:0] I_62,
  input [31:0] I_63,
  input [31:0] I_64,
  input [31:0] I_65,
  input [31:0] I_66,
  input [31:0] I_67,
  input [31:0] I_68,
  input [31:0] I_69,
  input [31:0] I_7,
  input [31:0] I_70,
  input [31:0] I_71,
  input [31:0] I_72,
  input [31:0] I_73,
  input [31:0] I_74,
  input [31:0] I_75,
  input [31:0] I_76,
  input [31:0] I_77,
  input [31:0] I_78,
  input [31:0] I_79,
  input [31:0] I_8,
  input [31:0] I_9,
  output [31:0] O,
  input [6:0] S
);


  wire [31:0] Mux80x32_inst0__I0;
  wire [31:0] Mux80x32_inst0__I1;
  wire [31:0] Mux80x32_inst0__I10;
  wire [31:0] Mux80x32_inst0__I11;
  wire [31:0] Mux80x32_inst0__I12;
  wire [31:0] Mux80x32_inst0__I13;
  wire [31:0] Mux80x32_inst0__I14;
  wire [31:0] Mux80x32_inst0__I15;
  wire [31:0] Mux80x32_inst0__I16;
  wire [31:0] Mux80x32_inst0__I17;
  wire [31:0] Mux80x32_inst0__I18;
  wire [31:0] Mux80x32_inst0__I19;
  wire [31:0] Mux80x32_inst0__I2;
  wire [31:0] Mux80x32_inst0__I20;
  wire [31:0] Mux80x32_inst0__I21;
  wire [31:0] Mux80x32_inst0__I22;
  wire [31:0] Mux80x32_inst0__I23;
  wire [31:0] Mux80x32_inst0__I24;
  wire [31:0] Mux80x32_inst0__I25;
  wire [31:0] Mux80x32_inst0__I26;
  wire [31:0] Mux80x32_inst0__I27;
  wire [31:0] Mux80x32_inst0__I28;
  wire [31:0] Mux80x32_inst0__I29;
  wire [31:0] Mux80x32_inst0__I3;
  wire [31:0] Mux80x32_inst0__I30;
  wire [31:0] Mux80x32_inst0__I31;
  wire [31:0] Mux80x32_inst0__I32;
  wire [31:0] Mux80x32_inst0__I33;
  wire [31:0] Mux80x32_inst0__I34;
  wire [31:0] Mux80x32_inst0__I35;
  wire [31:0] Mux80x32_inst0__I36;
  wire [31:0] Mux80x32_inst0__I37;
  wire [31:0] Mux80x32_inst0__I38;
  wire [31:0] Mux80x32_inst0__I39;
  wire [31:0] Mux80x32_inst0__I4;
  wire [31:0] Mux80x32_inst0__I40;
  wire [31:0] Mux80x32_inst0__I41;
  wire [31:0] Mux80x32_inst0__I42;
  wire [31:0] Mux80x32_inst0__I43;
  wire [31:0] Mux80x32_inst0__I44;
  wire [31:0] Mux80x32_inst0__I45;
  wire [31:0] Mux80x32_inst0__I46;
  wire [31:0] Mux80x32_inst0__I47;
  wire [31:0] Mux80x32_inst0__I48;
  wire [31:0] Mux80x32_inst0__I49;
  wire [31:0] Mux80x32_inst0__I5;
  wire [31:0] Mux80x32_inst0__I50;
  wire [31:0] Mux80x32_inst0__I51;
  wire [31:0] Mux80x32_inst0__I52;
  wire [31:0] Mux80x32_inst0__I53;
  wire [31:0] Mux80x32_inst0__I54;
  wire [31:0] Mux80x32_inst0__I55;
  wire [31:0] Mux80x32_inst0__I56;
  wire [31:0] Mux80x32_inst0__I57;
  wire [31:0] Mux80x32_inst0__I58;
  wire [31:0] Mux80x32_inst0__I59;
  wire [31:0] Mux80x32_inst0__I6;
  wire [31:0] Mux80x32_inst0__I60;
  wire [31:0] Mux80x32_inst0__I61;
  wire [31:0] Mux80x32_inst0__I62;
  wire [31:0] Mux80x32_inst0__I63;
  wire [31:0] Mux80x32_inst0__I64;
  wire [31:0] Mux80x32_inst0__I65;
  wire [31:0] Mux80x32_inst0__I66;
  wire [31:0] Mux80x32_inst0__I67;
  wire [31:0] Mux80x32_inst0__I68;
  wire [31:0] Mux80x32_inst0__I69;
  wire [31:0] Mux80x32_inst0__I7;
  wire [31:0] Mux80x32_inst0__I70;
  wire [31:0] Mux80x32_inst0__I71;
  wire [31:0] Mux80x32_inst0__I72;
  wire [31:0] Mux80x32_inst0__I73;
  wire [31:0] Mux80x32_inst0__I74;
  wire [31:0] Mux80x32_inst0__I75;
  wire [31:0] Mux80x32_inst0__I76;
  wire [31:0] Mux80x32_inst0__I77;
  wire [31:0] Mux80x32_inst0__I78;
  wire [31:0] Mux80x32_inst0__I79;
  wire [31:0] Mux80x32_inst0__I8;
  wire [31:0] Mux80x32_inst0__I9;
  wire [31:0] Mux80x32_inst0__O;
  wire [6:0] Mux80x32_inst0__S;
  Mux80x32 Mux80x32_inst0(
    .I0(Mux80x32_inst0__I0),
    .I1(Mux80x32_inst0__I1),
    .I10(Mux80x32_inst0__I10),
    .I11(Mux80x32_inst0__I11),
    .I12(Mux80x32_inst0__I12),
    .I13(Mux80x32_inst0__I13),
    .I14(Mux80x32_inst0__I14),
    .I15(Mux80x32_inst0__I15),
    .I16(Mux80x32_inst0__I16),
    .I17(Mux80x32_inst0__I17),
    .I18(Mux80x32_inst0__I18),
    .I19(Mux80x32_inst0__I19),
    .I2(Mux80x32_inst0__I2),
    .I20(Mux80x32_inst0__I20),
    .I21(Mux80x32_inst0__I21),
    .I22(Mux80x32_inst0__I22),
    .I23(Mux80x32_inst0__I23),
    .I24(Mux80x32_inst0__I24),
    .I25(Mux80x32_inst0__I25),
    .I26(Mux80x32_inst0__I26),
    .I27(Mux80x32_inst0__I27),
    .I28(Mux80x32_inst0__I28),
    .I29(Mux80x32_inst0__I29),
    .I3(Mux80x32_inst0__I3),
    .I30(Mux80x32_inst0__I30),
    .I31(Mux80x32_inst0__I31),
    .I32(Mux80x32_inst0__I32),
    .I33(Mux80x32_inst0__I33),
    .I34(Mux80x32_inst0__I34),
    .I35(Mux80x32_inst0__I35),
    .I36(Mux80x32_inst0__I36),
    .I37(Mux80x32_inst0__I37),
    .I38(Mux80x32_inst0__I38),
    .I39(Mux80x32_inst0__I39),
    .I4(Mux80x32_inst0__I4),
    .I40(Mux80x32_inst0__I40),
    .I41(Mux80x32_inst0__I41),
    .I42(Mux80x32_inst0__I42),
    .I43(Mux80x32_inst0__I43),
    .I44(Mux80x32_inst0__I44),
    .I45(Mux80x32_inst0__I45),
    .I46(Mux80x32_inst0__I46),
    .I47(Mux80x32_inst0__I47),
    .I48(Mux80x32_inst0__I48),
    .I49(Mux80x32_inst0__I49),
    .I5(Mux80x32_inst0__I5),
    .I50(Mux80x32_inst0__I50),
    .I51(Mux80x32_inst0__I51),
    .I52(Mux80x32_inst0__I52),
    .I53(Mux80x32_inst0__I53),
    .I54(Mux80x32_inst0__I54),
    .I55(Mux80x32_inst0__I55),
    .I56(Mux80x32_inst0__I56),
    .I57(Mux80x32_inst0__I57),
    .I58(Mux80x32_inst0__I58),
    .I59(Mux80x32_inst0__I59),
    .I6(Mux80x32_inst0__I6),
    .I60(Mux80x32_inst0__I60),
    .I61(Mux80x32_inst0__I61),
    .I62(Mux80x32_inst0__I62),
    .I63(Mux80x32_inst0__I63),
    .I64(Mux80x32_inst0__I64),
    .I65(Mux80x32_inst0__I65),
    .I66(Mux80x32_inst0__I66),
    .I67(Mux80x32_inst0__I67),
    .I68(Mux80x32_inst0__I68),
    .I69(Mux80x32_inst0__I69),
    .I7(Mux80x32_inst0__I7),
    .I70(Mux80x32_inst0__I70),
    .I71(Mux80x32_inst0__I71),
    .I72(Mux80x32_inst0__I72),
    .I73(Mux80x32_inst0__I73),
    .I74(Mux80x32_inst0__I74),
    .I75(Mux80x32_inst0__I75),
    .I76(Mux80x32_inst0__I76),
    .I77(Mux80x32_inst0__I77),
    .I78(Mux80x32_inst0__I78),
    .I79(Mux80x32_inst0__I79),
    .I8(Mux80x32_inst0__I8),
    .I9(Mux80x32_inst0__I9),
    .O(Mux80x32_inst0__O),
    .S(Mux80x32_inst0__S)
  );

  assign Mux80x32_inst0__I0[31:0] = I_0[31:0];

  assign Mux80x32_inst0__I1[31:0] = I_1[31:0];

  assign Mux80x32_inst0__I10[31:0] = I_10[31:0];

  assign Mux80x32_inst0__I11[31:0] = I_11[31:0];

  assign Mux80x32_inst0__I12[31:0] = I_12[31:0];

  assign Mux80x32_inst0__I13[31:0] = I_13[31:0];

  assign Mux80x32_inst0__I14[31:0] = I_14[31:0];

  assign Mux80x32_inst0__I15[31:0] = I_15[31:0];

  assign Mux80x32_inst0__I16[31:0] = I_16[31:0];

  assign Mux80x32_inst0__I17[31:0] = I_17[31:0];

  assign Mux80x32_inst0__I18[31:0] = I_18[31:0];

  assign Mux80x32_inst0__I19[31:0] = I_19[31:0];

  assign Mux80x32_inst0__I2[31:0] = I_2[31:0];

  assign Mux80x32_inst0__I20[31:0] = I_20[31:0];

  assign Mux80x32_inst0__I21[31:0] = I_21[31:0];

  assign Mux80x32_inst0__I22[31:0] = I_22[31:0];

  assign Mux80x32_inst0__I23[31:0] = I_23[31:0];

  assign Mux80x32_inst0__I24[31:0] = I_24[31:0];

  assign Mux80x32_inst0__I25[31:0] = I_25[31:0];

  assign Mux80x32_inst0__I26[31:0] = I_26[31:0];

  assign Mux80x32_inst0__I27[31:0] = I_27[31:0];

  assign Mux80x32_inst0__I28[31:0] = I_28[31:0];

  assign Mux80x32_inst0__I29[31:0] = I_29[31:0];

  assign Mux80x32_inst0__I3[31:0] = I_3[31:0];

  assign Mux80x32_inst0__I30[31:0] = I_30[31:0];

  assign Mux80x32_inst0__I31[31:0] = I_31[31:0];

  assign Mux80x32_inst0__I32[31:0] = I_32[31:0];

  assign Mux80x32_inst0__I33[31:0] = I_33[31:0];

  assign Mux80x32_inst0__I34[31:0] = I_34[31:0];

  assign Mux80x32_inst0__I35[31:0] = I_35[31:0];

  assign Mux80x32_inst0__I36[31:0] = I_36[31:0];

  assign Mux80x32_inst0__I37[31:0] = I_37[31:0];

  assign Mux80x32_inst0__I38[31:0] = I_38[31:0];

  assign Mux80x32_inst0__I39[31:0] = I_39[31:0];

  assign Mux80x32_inst0__I4[31:0] = I_4[31:0];

  assign Mux80x32_inst0__I40[31:0] = I_40[31:0];

  assign Mux80x32_inst0__I41[31:0] = I_41[31:0];

  assign Mux80x32_inst0__I42[31:0] = I_42[31:0];

  assign Mux80x32_inst0__I43[31:0] = I_43[31:0];

  assign Mux80x32_inst0__I44[31:0] = I_44[31:0];

  assign Mux80x32_inst0__I45[31:0] = I_45[31:0];

  assign Mux80x32_inst0__I46[31:0] = I_46[31:0];

  assign Mux80x32_inst0__I47[31:0] = I_47[31:0];

  assign Mux80x32_inst0__I48[31:0] = I_48[31:0];

  assign Mux80x32_inst0__I49[31:0] = I_49[31:0];

  assign Mux80x32_inst0__I5[31:0] = I_5[31:0];

  assign Mux80x32_inst0__I50[31:0] = I_50[31:0];

  assign Mux80x32_inst0__I51[31:0] = I_51[31:0];

  assign Mux80x32_inst0__I52[31:0] = I_52[31:0];

  assign Mux80x32_inst0__I53[31:0] = I_53[31:0];

  assign Mux80x32_inst0__I54[31:0] = I_54[31:0];

  assign Mux80x32_inst0__I55[31:0] = I_55[31:0];

  assign Mux80x32_inst0__I56[31:0] = I_56[31:0];

  assign Mux80x32_inst0__I57[31:0] = I_57[31:0];

  assign Mux80x32_inst0__I58[31:0] = I_58[31:0];

  assign Mux80x32_inst0__I59[31:0] = I_59[31:0];

  assign Mux80x32_inst0__I6[31:0] = I_6[31:0];

  assign Mux80x32_inst0__I60[31:0] = I_60[31:0];

  assign Mux80x32_inst0__I61[31:0] = I_61[31:0];

  assign Mux80x32_inst0__I62[31:0] = I_62[31:0];

  assign Mux80x32_inst0__I63[31:0] = I_63[31:0];

  assign Mux80x32_inst0__I64[31:0] = I_64[31:0];

  assign Mux80x32_inst0__I65[31:0] = I_65[31:0];

  assign Mux80x32_inst0__I66[31:0] = I_66[31:0];

  assign Mux80x32_inst0__I67[31:0] = I_67[31:0];

  assign Mux80x32_inst0__I68[31:0] = I_68[31:0];

  assign Mux80x32_inst0__I69[31:0] = I_69[31:0];

  assign Mux80x32_inst0__I7[31:0] = I_7[31:0];

  assign Mux80x32_inst0__I70[31:0] = I_70[31:0];

  assign Mux80x32_inst0__I71[31:0] = I_71[31:0];

  assign Mux80x32_inst0__I72[31:0] = I_72[31:0];

  assign Mux80x32_inst0__I73[31:0] = I_73[31:0];

  assign Mux80x32_inst0__I74[31:0] = I_74[31:0];

  assign Mux80x32_inst0__I75[31:0] = I_75[31:0];

  assign Mux80x32_inst0__I76[31:0] = I_76[31:0];

  assign Mux80x32_inst0__I77[31:0] = I_77[31:0];

  assign Mux80x32_inst0__I78[31:0] = I_78[31:0];

  assign Mux80x32_inst0__I79[31:0] = I_79[31:0];

  assign Mux80x32_inst0__I8[31:0] = I_8[31:0];

  assign Mux80x32_inst0__I9[31:0] = I_9[31:0];

  assign O[31:0] = Mux80x32_inst0__O[31:0];

  assign Mux80x32_inst0__S[6:0] = S[6:0];


endmodule  // MuxWrapper_80_32

module Mux7x32 (
  input [31:0] I0,
  input [31:0] I1,
  input [31:0] I2,
  input [31:0] I3,
  input [31:0] I4,
  input [31:0] I5,
  input [31:0] I6,
  output [31:0] O,
  input [2:0] S
);


  // Instancing generated Module: commonlib.muxn(N:7, width:32)
  wire [31:0] coreir_commonlib_mux7x32_inst0__in_data_0;
  wire [31:0] coreir_commonlib_mux7x32_inst0__in_data_1;
  wire [31:0] coreir_commonlib_mux7x32_inst0__in_data_2;
  wire [31:0] coreir_commonlib_mux7x32_inst0__in_data_3;
  wire [31:0] coreir_commonlib_mux7x32_inst0__in_data_4;
  wire [31:0] coreir_commonlib_mux7x32_inst0__in_data_5;
  wire [31:0] coreir_commonlib_mux7x32_inst0__in_data_6;
  wire [2:0] coreir_commonlib_mux7x32_inst0__in_sel;
  wire [31:0] coreir_commonlib_mux7x32_inst0__out;
  commonlib_muxn__N7__width32 coreir_commonlib_mux7x32_inst0(
    .in_data_0(coreir_commonlib_mux7x32_inst0__in_data_0),
    .in_data_1(coreir_commonlib_mux7x32_inst0__in_data_1),
    .in_data_2(coreir_commonlib_mux7x32_inst0__in_data_2),
    .in_data_3(coreir_commonlib_mux7x32_inst0__in_data_3),
    .in_data_4(coreir_commonlib_mux7x32_inst0__in_data_4),
    .in_data_5(coreir_commonlib_mux7x32_inst0__in_data_5),
    .in_data_6(coreir_commonlib_mux7x32_inst0__in_data_6),
    .in_sel(coreir_commonlib_mux7x32_inst0__in_sel),
    .out(coreir_commonlib_mux7x32_inst0__out)
  );

  assign coreir_commonlib_mux7x32_inst0__in_data_0[31:0] = I0[31:0];

  assign coreir_commonlib_mux7x32_inst0__in_data_1[31:0] = I1[31:0];

  assign coreir_commonlib_mux7x32_inst0__in_data_2[31:0] = I2[31:0];

  assign coreir_commonlib_mux7x32_inst0__in_data_3[31:0] = I3[31:0];

  assign coreir_commonlib_mux7x32_inst0__in_data_4[31:0] = I4[31:0];

  assign coreir_commonlib_mux7x32_inst0__in_data_5[31:0] = I5[31:0];

  assign coreir_commonlib_mux7x32_inst0__in_data_6[31:0] = I6[31:0];

  assign coreir_commonlib_mux7x32_inst0__in_sel[2:0] = S[2:0];

  assign O[31:0] = coreir_commonlib_mux7x32_inst0__out[31:0];


endmodule  // Mux7x32

module MuxWrapper_7_32 (
  input [31:0] I_0,
  input [31:0] I_1,
  input [31:0] I_2,
  input [31:0] I_3,
  input [31:0] I_4,
  input [31:0] I_5,
  input [31:0] I_6,
  output [31:0] O,
  input [2:0] S
);


  wire [31:0] Mux7x32_inst0__I0;
  wire [31:0] Mux7x32_inst0__I1;
  wire [31:0] Mux7x32_inst0__I2;
  wire [31:0] Mux7x32_inst0__I3;
  wire [31:0] Mux7x32_inst0__I4;
  wire [31:0] Mux7x32_inst0__I5;
  wire [31:0] Mux7x32_inst0__I6;
  wire [31:0] Mux7x32_inst0__O;
  wire [2:0] Mux7x32_inst0__S;
  Mux7x32 Mux7x32_inst0(
    .I0(Mux7x32_inst0__I0),
    .I1(Mux7x32_inst0__I1),
    .I2(Mux7x32_inst0__I2),
    .I3(Mux7x32_inst0__I3),
    .I4(Mux7x32_inst0__I4),
    .I5(Mux7x32_inst0__I5),
    .I6(Mux7x32_inst0__I6),
    .O(Mux7x32_inst0__O),
    .S(Mux7x32_inst0__S)
  );

  assign Mux7x32_inst0__I0[31:0] = I_0[31:0];

  assign Mux7x32_inst0__I1[31:0] = I_1[31:0];

  assign Mux7x32_inst0__I2[31:0] = I_2[31:0];

  assign Mux7x32_inst0__I3[31:0] = I_3[31:0];

  assign Mux7x32_inst0__I4[31:0] = I_4[31:0];

  assign Mux7x32_inst0__I5[31:0] = I_5[31:0];

  assign Mux7x32_inst0__I6[31:0] = I_6[31:0];

  assign O[31:0] = Mux7x32_inst0__O[31:0];

  assign Mux7x32_inst0__S[2:0] = S[2:0];


endmodule  // MuxWrapper_7_32

module Mux4x16 (
  input [15:0] I0,
  input [15:0] I1,
  input [15:0] I2,
  input [15:0] I3,
  output [15:0] O,
  input [1:0] S
);


  // Instancing generated Module: commonlib.muxn(N:4, width:16)
  wire [15:0] coreir_commonlib_mux4x16_inst0__in_data_0;
  wire [15:0] coreir_commonlib_mux4x16_inst0__in_data_1;
  wire [15:0] coreir_commonlib_mux4x16_inst0__in_data_2;
  wire [15:0] coreir_commonlib_mux4x16_inst0__in_data_3;
  wire [1:0] coreir_commonlib_mux4x16_inst0__in_sel;
  wire [15:0] coreir_commonlib_mux4x16_inst0__out;
  commonlib_muxn__N4__width16 coreir_commonlib_mux4x16_inst0(
    .in_data_0(coreir_commonlib_mux4x16_inst0__in_data_0),
    .in_data_1(coreir_commonlib_mux4x16_inst0__in_data_1),
    .in_data_2(coreir_commonlib_mux4x16_inst0__in_data_2),
    .in_data_3(coreir_commonlib_mux4x16_inst0__in_data_3),
    .in_sel(coreir_commonlib_mux4x16_inst0__in_sel),
    .out(coreir_commonlib_mux4x16_inst0__out)
  );

  assign coreir_commonlib_mux4x16_inst0__in_data_0[15:0] = I0[15:0];

  assign coreir_commonlib_mux4x16_inst0__in_data_1[15:0] = I1[15:0];

  assign coreir_commonlib_mux4x16_inst0__in_data_2[15:0] = I2[15:0];

  assign coreir_commonlib_mux4x16_inst0__in_data_3[15:0] = I3[15:0];

  assign coreir_commonlib_mux4x16_inst0__in_sel[1:0] = S[1:0];

  assign O[15:0] = coreir_commonlib_mux4x16_inst0__out[15:0];


endmodule  // Mux4x16

module MuxWrapper_4_16 (
  input [15:0] I_0,
  input [15:0] I_1,
  input [15:0] I_2,
  input [15:0] I_3,
  output [15:0] O,
  input [1:0] S
);


  wire [15:0] Mux4x16_inst0__I0;
  wire [15:0] Mux4x16_inst0__I1;
  wire [15:0] Mux4x16_inst0__I2;
  wire [15:0] Mux4x16_inst0__I3;
  wire [15:0] Mux4x16_inst0__O;
  wire [1:0] Mux4x16_inst0__S;
  Mux4x16 Mux4x16_inst0(
    .I0(Mux4x16_inst0__I0),
    .I1(Mux4x16_inst0__I1),
    .I2(Mux4x16_inst0__I2),
    .I3(Mux4x16_inst0__I3),
    .O(Mux4x16_inst0__O),
    .S(Mux4x16_inst0__S)
  );

  assign Mux4x16_inst0__I0[15:0] = I_0[15:0];

  assign Mux4x16_inst0__I1[15:0] = I_1[15:0];

  assign Mux4x16_inst0__I2[15:0] = I_2[15:0];

  assign Mux4x16_inst0__I3[15:0] = I_3[15:0];

  assign O[15:0] = Mux4x16_inst0__O[15:0];

  assign Mux4x16_inst0__S[1:0] = S[1:0];


endmodule  // MuxWrapper_4_16

module Mux4x1 (
  input [0:0] I0,
  input [0:0] I1,
  input [0:0] I2,
  input [0:0] I3,
  output [0:0] O,
  input [1:0] S
);


  // Instancing generated Module: commonlib.muxn(N:4, width:1)
  wire [0:0] coreir_commonlib_mux4x1_inst0__in_data_0;
  wire [0:0] coreir_commonlib_mux4x1_inst0__in_data_1;
  wire [0:0] coreir_commonlib_mux4x1_inst0__in_data_2;
  wire [0:0] coreir_commonlib_mux4x1_inst0__in_data_3;
  wire [1:0] coreir_commonlib_mux4x1_inst0__in_sel;
  wire [0:0] coreir_commonlib_mux4x1_inst0__out;
  commonlib_muxn__N4__width1 coreir_commonlib_mux4x1_inst0(
    .in_data_0(coreir_commonlib_mux4x1_inst0__in_data_0),
    .in_data_1(coreir_commonlib_mux4x1_inst0__in_data_1),
    .in_data_2(coreir_commonlib_mux4x1_inst0__in_data_2),
    .in_data_3(coreir_commonlib_mux4x1_inst0__in_data_3),
    .in_sel(coreir_commonlib_mux4x1_inst0__in_sel),
    .out(coreir_commonlib_mux4x1_inst0__out)
  );

  assign coreir_commonlib_mux4x1_inst0__in_data_0[0:0] = I0[0:0];

  assign coreir_commonlib_mux4x1_inst0__in_data_1[0:0] = I1[0:0];

  assign coreir_commonlib_mux4x1_inst0__in_data_2[0:0] = I2[0:0];

  assign coreir_commonlib_mux4x1_inst0__in_data_3[0:0] = I3[0:0];

  assign coreir_commonlib_mux4x1_inst0__in_sel[1:0] = S[1:0];

  assign O[0:0] = coreir_commonlib_mux4x1_inst0__out[0:0];


endmodule  // Mux4x1

module MuxWrapper_4_1 (
  input [0:0] I_0,
  input [0:0] I_1,
  input [0:0] I_2,
  input [0:0] I_3,
  output [0:0] O,
  input [1:0] S
);


  wire [0:0] Mux4x1_inst0__I0;
  wire [0:0] Mux4x1_inst0__I1;
  wire [0:0] Mux4x1_inst0__I2;
  wire [0:0] Mux4x1_inst0__I3;
  wire [0:0] Mux4x1_inst0__O;
  wire [1:0] Mux4x1_inst0__S;
  Mux4x1 Mux4x1_inst0(
    .I0(Mux4x1_inst0__I0),
    .I1(Mux4x1_inst0__I1),
    .I2(Mux4x1_inst0__I2),
    .I3(Mux4x1_inst0__I3),
    .O(Mux4x1_inst0__O),
    .S(Mux4x1_inst0__S)
  );

  assign Mux4x1_inst0__I0[0:0] = I_0[0:0];

  assign Mux4x1_inst0__I1[0:0] = I_1[0:0];

  assign Mux4x1_inst0__I2[0:0] = I_2[0:0];

  assign Mux4x1_inst0__I3[0:0] = I_3[0:0];

  assign O[0:0] = Mux4x1_inst0__O[0:0];

  assign Mux4x1_inst0__S[1:0] = S[1:0];


endmodule  // MuxWrapper_4_1

module Mux2xOutBits4 (
  input [3:0] I0,
  input [3:0] I1,
  output [3:0] O,
  input  S
);


  // Instancing generated Module: commonlib.muxn(N:2, width:4)
  wire [3:0] coreir_commonlib_mux2x4_inst0__in_data_0;
  wire [3:0] coreir_commonlib_mux2x4_inst0__in_data_1;
  wire [0:0] coreir_commonlib_mux2x4_inst0__in_sel;
  wire [3:0] coreir_commonlib_mux2x4_inst0__out;
  commonlib_muxn__N2__width4 coreir_commonlib_mux2x4_inst0(
    .in_data_0(coreir_commonlib_mux2x4_inst0__in_data_0),
    .in_data_1(coreir_commonlib_mux2x4_inst0__in_data_1),
    .in_sel(coreir_commonlib_mux2x4_inst0__in_sel),
    .out(coreir_commonlib_mux2x4_inst0__out)
  );

  assign coreir_commonlib_mux2x4_inst0__in_data_0[3:0] = I0[3:0];

  assign coreir_commonlib_mux2x4_inst0__in_data_1[3:0] = I1[3:0];

  assign coreir_commonlib_mux2x4_inst0__in_sel[0] = S;

  assign O[3:0] = coreir_commonlib_mux2x4_inst0__out[3:0];


endmodule  // Mux2xOutBits4

module Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_4 (
  input  ASYNCRESET,
  input  CE,
  input  CLK,
  input [3:0] I,
  output [3:0] O
);


  wire [3:0] enable_mux__I0;
  wire [3:0] enable_mux__I1;
  wire [3:0] enable_mux__O;
  wire  enable_mux__S;
  Mux2xOutBits4 enable_mux(
    .I0(enable_mux__I0),
    .I1(enable_mux__I1),
    .O(enable_mux__O),
    .S(enable_mux__S)
  );

  // Instancing generated Module: coreir.reg_arst(width:4)
  wire  value__arst;
  wire  value__clk;
  wire [3:0] value__in;
  wire [3:0] value__out;
  coreir_reg_arst #(.arst_posedge(1),.clk_posedge(1),.init(4'h0),.width(4)) value(
    .arst(value__arst),
    .clk(value__clk),
    .in(value__in),
    .out(value__out)
  );

  assign enable_mux__I0[3:0] = value__out[3:0];

  assign enable_mux__I1[3:0] = I[3:0];

  assign value__in[3:0] = enable_mux__O[3:0];

  assign enable_mux__S = CE;

  assign value__arst = ASYNCRESET;

  assign value__clk = CLK;

  assign O[3:0] = value__out[3:0];


endmodule  // Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_4

module Mux2xOutBits2 (
  input [1:0] I0,
  input [1:0] I1,
  output [1:0] O,
  input  S
);


  // Instancing generated Module: commonlib.muxn(N:2, width:2)
  wire [1:0] coreir_commonlib_mux2x2_inst0__in_data_0;
  wire [1:0] coreir_commonlib_mux2x2_inst0__in_data_1;
  wire [0:0] coreir_commonlib_mux2x2_inst0__in_sel;
  wire [1:0] coreir_commonlib_mux2x2_inst0__out;
  commonlib_muxn__N2__width2 coreir_commonlib_mux2x2_inst0(
    .in_data_0(coreir_commonlib_mux2x2_inst0__in_data_0),
    .in_data_1(coreir_commonlib_mux2x2_inst0__in_data_1),
    .in_sel(coreir_commonlib_mux2x2_inst0__in_sel),
    .out(coreir_commonlib_mux2x2_inst0__out)
  );

  assign coreir_commonlib_mux2x2_inst0__in_data_0[1:0] = I0[1:0];

  assign coreir_commonlib_mux2x2_inst0__in_data_1[1:0] = I1[1:0];

  assign coreir_commonlib_mux2x2_inst0__in_sel[0] = S;

  assign O[1:0] = coreir_commonlib_mux2x2_inst0__out[1:0];


endmodule  // Mux2xOutBits2

module Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2 (
  input  ASYNCRESET,
  input  CE,
  input  CLK,
  input [1:0] I,
  output [1:0] O
);


  wire [1:0] enable_mux__I0;
  wire [1:0] enable_mux__I1;
  wire [1:0] enable_mux__O;
  wire  enable_mux__S;
  Mux2xOutBits2 enable_mux(
    .I0(enable_mux__I0),
    .I1(enable_mux__I1),
    .O(enable_mux__O),
    .S(enable_mux__S)
  );

  // Instancing generated Module: coreir.reg_arst(width:2)
  wire  value__arst;
  wire  value__clk;
  wire [1:0] value__in;
  wire [1:0] value__out;
  coreir_reg_arst #(.arst_posedge(1),.clk_posedge(1),.init(2'h0),.width(2)) value(
    .arst(value__arst),
    .clk(value__clk),
    .in(value__in),
    .out(value__out)
  );

  assign enable_mux__I0[1:0] = value__out[1:0];

  assign enable_mux__I1[1:0] = I[1:0];

  assign value__in[1:0] = enable_mux__O[1:0];

  assign enable_mux__S = CE;

  assign value__arst = ASYNCRESET;

  assign value__clk = CLK;

  assign O[1:0] = value__out[1:0];


endmodule  // Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2

module Mux2xOutBits1 (
  input [0:0] I0,
  input [0:0] I1,
  output [0:0] O,
  input  S
);


  // Instancing generated Module: commonlib.muxn(N:2, width:1)
  wire [0:0] coreir_commonlib_mux2x1_inst0__in_data_0;
  wire [0:0] coreir_commonlib_mux2x1_inst0__in_data_1;
  wire [0:0] coreir_commonlib_mux2x1_inst0__in_sel;
  wire [0:0] coreir_commonlib_mux2x1_inst0__out;
  commonlib_muxn__N2__width1 coreir_commonlib_mux2x1_inst0(
    .in_data_0(coreir_commonlib_mux2x1_inst0__in_data_0),
    .in_data_1(coreir_commonlib_mux2x1_inst0__in_data_1),
    .in_sel(coreir_commonlib_mux2x1_inst0__in_sel),
    .out(coreir_commonlib_mux2x1_inst0__out)
  );

  assign coreir_commonlib_mux2x1_inst0__in_data_0[0:0] = I0[0:0];

  assign coreir_commonlib_mux2x1_inst0__in_data_1[0:0] = I1[0:0];

  assign coreir_commonlib_mux2x1_inst0__in_sel[0] = S;

  assign O[0:0] = coreir_commonlib_mux2x1_inst0__out[0:0];


endmodule  // Mux2xOutBits1

module Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1 (
  input  ASYNCRESET,
  input  CE,
  input  CLK,
  input [0:0] I,
  output [0:0] O
);


  wire [0:0] enable_mux__I0;
  wire [0:0] enable_mux__I1;
  wire [0:0] enable_mux__O;
  wire  enable_mux__S;
  Mux2xOutBits1 enable_mux(
    .I0(enable_mux__I0),
    .I1(enable_mux__I1),
    .O(enable_mux__O),
    .S(enable_mux__S)
  );

  // Instancing generated Module: coreir.reg_arst(width:1)
  wire  value__arst;
  wire  value__clk;
  wire [0:0] value__in;
  wire [0:0] value__out;
  coreir_reg_arst #(.arst_posedge(1),.clk_posedge(1),.init(1'h0),.width(1)) value(
    .arst(value__arst),
    .clk(value__clk),
    .in(value__in),
    .out(value__out)
  );

  assign enable_mux__I0[0:0] = value__out[0:0];

  assign enable_mux__I1[0:0] = I[0:0];

  assign value__in[0:0] = enable_mux__O[0:0];

  assign enable_mux__S = CE;

  assign value__arst = ASYNCRESET;

  assign value__clk = CLK;

  assign O[0:0] = value__out[0:0];


endmodule  // Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1

module Mux2x32 (
  input [31:0] I0,
  input [31:0] I1,
  output [31:0] O,
  input  S
);


  // Instancing generated Module: commonlib.muxn(N:2, width:32)
  wire [31:0] coreir_commonlib_mux2x32_inst0__in_data_0;
  wire [31:0] coreir_commonlib_mux2x32_inst0__in_data_1;
  wire [0:0] coreir_commonlib_mux2x32_inst0__in_sel;
  wire [31:0] coreir_commonlib_mux2x32_inst0__out;
  commonlib_muxn__N2__width32 coreir_commonlib_mux2x32_inst0(
    .in_data_0(coreir_commonlib_mux2x32_inst0__in_data_0),
    .in_data_1(coreir_commonlib_mux2x32_inst0__in_data_1),
    .in_sel(coreir_commonlib_mux2x32_inst0__in_sel),
    .out(coreir_commonlib_mux2x32_inst0__out)
  );

  assign coreir_commonlib_mux2x32_inst0__in_data_0[31:0] = I0[31:0];

  assign coreir_commonlib_mux2x32_inst0__in_data_1[31:0] = I1[31:0];

  assign coreir_commonlib_mux2x32_inst0__in_sel[0] = S;

  assign O[31:0] = coreir_commonlib_mux2x32_inst0__out[31:0];


endmodule  // Mux2x32

module MuxWrapper_2_32 (
  input [31:0] I_0,
  input [31:0] I_1,
  output [31:0] O,
  input [0:0] S
);


  wire [31:0] Mux2x32_inst0__I0;
  wire [31:0] Mux2x32_inst0__I1;
  wire [31:0] Mux2x32_inst0__O;
  wire  Mux2x32_inst0__S;
  Mux2x32 Mux2x32_inst0(
    .I0(Mux2x32_inst0__I0),
    .I1(Mux2x32_inst0__I1),
    .O(Mux2x32_inst0__O),
    .S(Mux2x32_inst0__S)
  );

  assign Mux2x32_inst0__I0[31:0] = I_0[31:0];

  assign Mux2x32_inst0__I1[31:0] = I_1[31:0];

  assign O[31:0] = Mux2x32_inst0__O[31:0];

  assign Mux2x32_inst0__S = S[0];


endmodule  // MuxWrapper_2_32

module MuxWithDefaultWrapper_7_32_8_0 (
  input [0:0] EN,
  input [31:0] I_0,
  input [31:0] I_1,
  input [31:0] I_2,
  input [31:0] I_3,
  input [31:0] I_4,
  input [31:0] I_5,
  input [31:0] I_6,
  output [31:0] O,
  input [7:0] S
);


  wire [31:0] MuxWrapper_2_32_inst0__I_0;
  wire [31:0] MuxWrapper_2_32_inst0__I_1;
  wire [31:0] MuxWrapper_2_32_inst0__O;
  wire [0:0] MuxWrapper_2_32_inst0__S;
  MuxWrapper_2_32 MuxWrapper_2_32_inst0(
    .I_0(MuxWrapper_2_32_inst0__I_0),
    .I_1(MuxWrapper_2_32_inst0__I_1),
    .O(MuxWrapper_2_32_inst0__O),
    .S(MuxWrapper_2_32_inst0__S)
  );

  wire [31:0] MuxWrapper_7_32_inst0__I_0;
  wire [31:0] MuxWrapper_7_32_inst0__I_1;
  wire [31:0] MuxWrapper_7_32_inst0__I_2;
  wire [31:0] MuxWrapper_7_32_inst0__I_3;
  wire [31:0] MuxWrapper_7_32_inst0__I_4;
  wire [31:0] MuxWrapper_7_32_inst0__I_5;
  wire [31:0] MuxWrapper_7_32_inst0__I_6;
  wire [31:0] MuxWrapper_7_32_inst0__O;
  wire [2:0] MuxWrapper_7_32_inst0__S;
  MuxWrapper_7_32 MuxWrapper_7_32_inst0(
    .I_0(MuxWrapper_7_32_inst0__I_0),
    .I_1(MuxWrapper_7_32_inst0__I_1),
    .I_2(MuxWrapper_7_32_inst0__I_2),
    .I_3(MuxWrapper_7_32_inst0__I_3),
    .I_4(MuxWrapper_7_32_inst0__I_4),
    .I_5(MuxWrapper_7_32_inst0__I_5),
    .I_6(MuxWrapper_7_32_inst0__I_6),
    .O(MuxWrapper_7_32_inst0__O),
    .S(MuxWrapper_7_32_inst0__S)
  );

  wire  and_inst0__in0;
  wire  and_inst0__in1;
  wire  and_inst0__out;
  corebit_and and_inst0(
    .in0(and_inst0__in0),
    .in1(and_inst0__in1),
    .out(and_inst0__out)
  );

  // Instancing generated Module: coreir.const(width:32)
  wire [31:0] const_0_32__out;
  coreir_const #(.value(32'h00000000),.width(32)) const_0_32(
    .out(const_0_32__out)
  );

  // Instancing generated Module: coreir.const(width:8)
  wire [7:0] const_7_8__out;
  coreir_const #(.value(8'h07),.width(8)) const_7_8(
    .out(const_7_8__out)
  );

  // Instancing generated Module: coreir.ult(width:8)
  wire [7:0] coreir_ult8_inst0__in0;
  wire [7:0] coreir_ult8_inst0__in1;
  wire  coreir_ult8_inst0__out;
  coreir_ult #(.width(8)) coreir_ult8_inst0(
    .in0(coreir_ult8_inst0__in0),
    .in1(coreir_ult8_inst0__in1),
    .out(coreir_ult8_inst0__out)
  );

  assign MuxWrapper_2_32_inst0__I_0[31:0] = const_0_32__out[31:0];

  assign MuxWrapper_2_32_inst0__I_1[31:0] = MuxWrapper_7_32_inst0__O[31:0];

  assign O[31:0] = MuxWrapper_2_32_inst0__O[31:0];

  assign MuxWrapper_2_32_inst0__S[0] = and_inst0__out;

  assign MuxWrapper_7_32_inst0__I_0[31:0] = I_0[31:0];

  assign MuxWrapper_7_32_inst0__I_1[31:0] = I_1[31:0];

  assign MuxWrapper_7_32_inst0__I_2[31:0] = I_2[31:0];

  assign MuxWrapper_7_32_inst0__I_3[31:0] = I_3[31:0];

  assign MuxWrapper_7_32_inst0__I_4[31:0] = I_4[31:0];

  assign MuxWrapper_7_32_inst0__I_5[31:0] = I_5[31:0];

  assign MuxWrapper_7_32_inst0__I_6[31:0] = I_6[31:0];

  assign MuxWrapper_7_32_inst0__S[0] = S[0];

  assign MuxWrapper_7_32_inst0__S[1] = S[1];

  assign MuxWrapper_7_32_inst0__S[2] = S[2];

  assign and_inst0__in0 = coreir_ult8_inst0__out;

  assign and_inst0__in1 = EN[0];

  assign coreir_ult8_inst0__in1[7:0] = const_7_8__out[7:0];

  assign coreir_ult8_inst0__in0[7:0] = S[7:0];


endmodule  // MuxWithDefaultWrapper_7_32_8_0

module Mux2x16 (
  input [15:0] I0,
  input [15:0] I1,
  output [15:0] O,
  input  S
);


  // Instancing generated Module: commonlib.muxn(N:2, width:16)
  wire [15:0] coreir_commonlib_mux2x16_inst0__in_data_0;
  wire [15:0] coreir_commonlib_mux2x16_inst0__in_data_1;
  wire [0:0] coreir_commonlib_mux2x16_inst0__in_sel;
  wire [15:0] coreir_commonlib_mux2x16_inst0__out;
  commonlib_muxn__N2__width16 coreir_commonlib_mux2x16_inst0(
    .in_data_0(coreir_commonlib_mux2x16_inst0__in_data_0),
    .in_data_1(coreir_commonlib_mux2x16_inst0__in_data_1),
    .in_sel(coreir_commonlib_mux2x16_inst0__in_sel),
    .out(coreir_commonlib_mux2x16_inst0__out)
  );

  assign coreir_commonlib_mux2x16_inst0__in_data_0[15:0] = I0[15:0];

  assign coreir_commonlib_mux2x16_inst0__in_data_1[15:0] = I1[15:0];

  assign coreir_commonlib_mux2x16_inst0__in_sel[0] = S;

  assign O[15:0] = coreir_commonlib_mux2x16_inst0__out[15:0];


endmodule  // Mux2x16

module MuxWrapper_2_16 (
  input [15:0] I_0,
  input [15:0] I_1,
  output [15:0] O,
  input [0:0] S
);


  wire [15:0] Mux2x16_inst0__I0;
  wire [15:0] Mux2x16_inst0__I1;
  wire [15:0] Mux2x16_inst0__O;
  wire  Mux2x16_inst0__S;
  Mux2x16 Mux2x16_inst0(
    .I0(Mux2x16_inst0__I0),
    .I1(Mux2x16_inst0__I1),
    .O(Mux2x16_inst0__O),
    .S(Mux2x16_inst0__S)
  );

  assign Mux2x16_inst0__I0[15:0] = I_0[15:0];

  assign Mux2x16_inst0__I1[15:0] = I_1[15:0];

  assign O[15:0] = Mux2x16_inst0__O[15:0];

  assign Mux2x16_inst0__S = S[0];


endmodule  // MuxWrapper_2_16

module Mux2x1 (
  input [0:0] I0,
  input [0:0] I1,
  output [0:0] O,
  input  S
);


  // Instancing generated Module: commonlib.muxn(N:2, width:1)
  wire [0:0] coreir_commonlib_mux2x1_inst0__in_data_0;
  wire [0:0] coreir_commonlib_mux2x1_inst0__in_data_1;
  wire [0:0] coreir_commonlib_mux2x1_inst0__in_sel;
  wire [0:0] coreir_commonlib_mux2x1_inst0__out;
  commonlib_muxn__N2__width1 coreir_commonlib_mux2x1_inst0(
    .in_data_0(coreir_commonlib_mux2x1_inst0__in_data_0),
    .in_data_1(coreir_commonlib_mux2x1_inst0__in_data_1),
    .in_sel(coreir_commonlib_mux2x1_inst0__in_sel),
    .out(coreir_commonlib_mux2x1_inst0__out)
  );

  assign coreir_commonlib_mux2x1_inst0__in_data_0[0:0] = I0[0:0];

  assign coreir_commonlib_mux2x1_inst0__in_data_1[0:0] = I1[0:0];

  assign coreir_commonlib_mux2x1_inst0__in_sel[0] = S;

  assign O[0:0] = coreir_commonlib_mux2x1_inst0__out[0:0];


endmodule  // Mux2x1

module MuxWrapper_2_1 (
  input [0:0] I_0,
  input [0:0] I_1,
  output [0:0] O,
  input [0:0] S
);


  wire [0:0] Mux2x1_inst0__I0;
  wire [0:0] Mux2x1_inst0__I1;
  wire [0:0] Mux2x1_inst0__O;
  wire  Mux2x1_inst0__S;
  Mux2x1 Mux2x1_inst0(
    .I0(Mux2x1_inst0__I0),
    .I1(Mux2x1_inst0__I1),
    .O(Mux2x1_inst0__O),
    .S(Mux2x1_inst0__S)
  );

  assign Mux2x1_inst0__I0[0:0] = I_0[0:0];

  assign Mux2x1_inst0__I1[0:0] = I_1[0:0];

  assign O[0:0] = Mux2x1_inst0__O[0:0];

  assign Mux2x1_inst0__S = S[0];


endmodule  // MuxWrapper_2_1

module Mux10x16 (
  input [15:0] I0,
  input [15:0] I1,
  input [15:0] I2,
  input [15:0] I3,
  input [15:0] I4,
  input [15:0] I5,
  input [15:0] I6,
  input [15:0] I7,
  input [15:0] I8,
  input [15:0] I9,
  output [15:0] O,
  input [3:0] S
);


  // Instancing generated Module: commonlib.muxn(N:10, width:16)
  wire [15:0] coreir_commonlib_mux10x16_inst0__in_data_0;
  wire [15:0] coreir_commonlib_mux10x16_inst0__in_data_1;
  wire [15:0] coreir_commonlib_mux10x16_inst0__in_data_2;
  wire [15:0] coreir_commonlib_mux10x16_inst0__in_data_3;
  wire [15:0] coreir_commonlib_mux10x16_inst0__in_data_4;
  wire [15:0] coreir_commonlib_mux10x16_inst0__in_data_5;
  wire [15:0] coreir_commonlib_mux10x16_inst0__in_data_6;
  wire [15:0] coreir_commonlib_mux10x16_inst0__in_data_7;
  wire [15:0] coreir_commonlib_mux10x16_inst0__in_data_8;
  wire [15:0] coreir_commonlib_mux10x16_inst0__in_data_9;
  wire [3:0] coreir_commonlib_mux10x16_inst0__in_sel;
  wire [15:0] coreir_commonlib_mux10x16_inst0__out;
  commonlib_muxn__N10__width16 coreir_commonlib_mux10x16_inst0(
    .in_data_0(coreir_commonlib_mux10x16_inst0__in_data_0),
    .in_data_1(coreir_commonlib_mux10x16_inst0__in_data_1),
    .in_data_2(coreir_commonlib_mux10x16_inst0__in_data_2),
    .in_data_3(coreir_commonlib_mux10x16_inst0__in_data_3),
    .in_data_4(coreir_commonlib_mux10x16_inst0__in_data_4),
    .in_data_5(coreir_commonlib_mux10x16_inst0__in_data_5),
    .in_data_6(coreir_commonlib_mux10x16_inst0__in_data_6),
    .in_data_7(coreir_commonlib_mux10x16_inst0__in_data_7),
    .in_data_8(coreir_commonlib_mux10x16_inst0__in_data_8),
    .in_data_9(coreir_commonlib_mux10x16_inst0__in_data_9),
    .in_sel(coreir_commonlib_mux10x16_inst0__in_sel),
    .out(coreir_commonlib_mux10x16_inst0__out)
  );

  assign coreir_commonlib_mux10x16_inst0__in_data_0[15:0] = I0[15:0];

  assign coreir_commonlib_mux10x16_inst0__in_data_1[15:0] = I1[15:0];

  assign coreir_commonlib_mux10x16_inst0__in_data_2[15:0] = I2[15:0];

  assign coreir_commonlib_mux10x16_inst0__in_data_3[15:0] = I3[15:0];

  assign coreir_commonlib_mux10x16_inst0__in_data_4[15:0] = I4[15:0];

  assign coreir_commonlib_mux10x16_inst0__in_data_5[15:0] = I5[15:0];

  assign coreir_commonlib_mux10x16_inst0__in_data_6[15:0] = I6[15:0];

  assign coreir_commonlib_mux10x16_inst0__in_data_7[15:0] = I7[15:0];

  assign coreir_commonlib_mux10x16_inst0__in_data_8[15:0] = I8[15:0];

  assign coreir_commonlib_mux10x16_inst0__in_data_9[15:0] = I9[15:0];

  assign coreir_commonlib_mux10x16_inst0__in_sel[3:0] = S[3:0];

  assign O[15:0] = coreir_commonlib_mux10x16_inst0__out[15:0];


endmodule  // Mux10x16

module MuxWrapper_10_16 (
  input [15:0] I_0,
  input [15:0] I_1,
  input [15:0] I_2,
  input [15:0] I_3,
  input [15:0] I_4,
  input [15:0] I_5,
  input [15:0] I_6,
  input [15:0] I_7,
  input [15:0] I_8,
  input [15:0] I_9,
  output [15:0] O,
  input [3:0] S
);


  wire [15:0] Mux10x16_inst0__I0;
  wire [15:0] Mux10x16_inst0__I1;
  wire [15:0] Mux10x16_inst0__I2;
  wire [15:0] Mux10x16_inst0__I3;
  wire [15:0] Mux10x16_inst0__I4;
  wire [15:0] Mux10x16_inst0__I5;
  wire [15:0] Mux10x16_inst0__I6;
  wire [15:0] Mux10x16_inst0__I7;
  wire [15:0] Mux10x16_inst0__I8;
  wire [15:0] Mux10x16_inst0__I9;
  wire [15:0] Mux10x16_inst0__O;
  wire [3:0] Mux10x16_inst0__S;
  Mux10x16 Mux10x16_inst0(
    .I0(Mux10x16_inst0__I0),
    .I1(Mux10x16_inst0__I1),
    .I2(Mux10x16_inst0__I2),
    .I3(Mux10x16_inst0__I3),
    .I4(Mux10x16_inst0__I4),
    .I5(Mux10x16_inst0__I5),
    .I6(Mux10x16_inst0__I6),
    .I7(Mux10x16_inst0__I7),
    .I8(Mux10x16_inst0__I8),
    .I9(Mux10x16_inst0__I9),
    .O(Mux10x16_inst0__O),
    .S(Mux10x16_inst0__S)
  );

  assign Mux10x16_inst0__I0[15:0] = I_0[15:0];

  assign Mux10x16_inst0__I1[15:0] = I_1[15:0];

  assign Mux10x16_inst0__I2[15:0] = I_2[15:0];

  assign Mux10x16_inst0__I3[15:0] = I_3[15:0];

  assign Mux10x16_inst0__I4[15:0] = I_4[15:0];

  assign Mux10x16_inst0__I5[15:0] = I_5[15:0];

  assign Mux10x16_inst0__I6[15:0] = I_6[15:0];

  assign Mux10x16_inst0__I7[15:0] = I_7[15:0];

  assign Mux10x16_inst0__I8[15:0] = I_8[15:0];

  assign Mux10x16_inst0__I9[15:0] = I_9[15:0];

  assign O[15:0] = Mux10x16_inst0__O[15:0];

  assign Mux10x16_inst0__S[3:0] = S[3:0];


endmodule  // MuxWrapper_10_16

module Mux10x1 (
  input [0:0] I0,
  input [0:0] I1,
  input [0:0] I2,
  input [0:0] I3,
  input [0:0] I4,
  input [0:0] I5,
  input [0:0] I6,
  input [0:0] I7,
  input [0:0] I8,
  input [0:0] I9,
  output [0:0] O,
  input [3:0] S
);


  // Instancing generated Module: commonlib.muxn(N:10, width:1)
  wire [0:0] coreir_commonlib_mux10x1_inst0__in_data_0;
  wire [0:0] coreir_commonlib_mux10x1_inst0__in_data_1;
  wire [0:0] coreir_commonlib_mux10x1_inst0__in_data_2;
  wire [0:0] coreir_commonlib_mux10x1_inst0__in_data_3;
  wire [0:0] coreir_commonlib_mux10x1_inst0__in_data_4;
  wire [0:0] coreir_commonlib_mux10x1_inst0__in_data_5;
  wire [0:0] coreir_commonlib_mux10x1_inst0__in_data_6;
  wire [0:0] coreir_commonlib_mux10x1_inst0__in_data_7;
  wire [0:0] coreir_commonlib_mux10x1_inst0__in_data_8;
  wire [0:0] coreir_commonlib_mux10x1_inst0__in_data_9;
  wire [3:0] coreir_commonlib_mux10x1_inst0__in_sel;
  wire [0:0] coreir_commonlib_mux10x1_inst0__out;
  commonlib_muxn__N10__width1 coreir_commonlib_mux10x1_inst0(
    .in_data_0(coreir_commonlib_mux10x1_inst0__in_data_0),
    .in_data_1(coreir_commonlib_mux10x1_inst0__in_data_1),
    .in_data_2(coreir_commonlib_mux10x1_inst0__in_data_2),
    .in_data_3(coreir_commonlib_mux10x1_inst0__in_data_3),
    .in_data_4(coreir_commonlib_mux10x1_inst0__in_data_4),
    .in_data_5(coreir_commonlib_mux10x1_inst0__in_data_5),
    .in_data_6(coreir_commonlib_mux10x1_inst0__in_data_6),
    .in_data_7(coreir_commonlib_mux10x1_inst0__in_data_7),
    .in_data_8(coreir_commonlib_mux10x1_inst0__in_data_8),
    .in_data_9(coreir_commonlib_mux10x1_inst0__in_data_9),
    .in_sel(coreir_commonlib_mux10x1_inst0__in_sel),
    .out(coreir_commonlib_mux10x1_inst0__out)
  );

  assign coreir_commonlib_mux10x1_inst0__in_data_0[0:0] = I0[0:0];

  assign coreir_commonlib_mux10x1_inst0__in_data_1[0:0] = I1[0:0];

  assign coreir_commonlib_mux10x1_inst0__in_data_2[0:0] = I2[0:0];

  assign coreir_commonlib_mux10x1_inst0__in_data_3[0:0] = I3[0:0];

  assign coreir_commonlib_mux10x1_inst0__in_data_4[0:0] = I4[0:0];

  assign coreir_commonlib_mux10x1_inst0__in_data_5[0:0] = I5[0:0];

  assign coreir_commonlib_mux10x1_inst0__in_data_6[0:0] = I6[0:0];

  assign coreir_commonlib_mux10x1_inst0__in_data_7[0:0] = I7[0:0];

  assign coreir_commonlib_mux10x1_inst0__in_data_8[0:0] = I8[0:0];

  assign coreir_commonlib_mux10x1_inst0__in_data_9[0:0] = I9[0:0];

  assign coreir_commonlib_mux10x1_inst0__in_sel[3:0] = S[3:0];

  assign O[0:0] = coreir_commonlib_mux10x1_inst0__out[0:0];


endmodule  // Mux10x1

module MuxWrapper_10_1 (
  input [0:0] I_0,
  input [0:0] I_1,
  input [0:0] I_2,
  input [0:0] I_3,
  input [0:0] I_4,
  input [0:0] I_5,
  input [0:0] I_6,
  input [0:0] I_7,
  input [0:0] I_8,
  input [0:0] I_9,
  output [0:0] O,
  input [3:0] S
);


  wire [0:0] Mux10x1_inst0__I0;
  wire [0:0] Mux10x1_inst0__I1;
  wire [0:0] Mux10x1_inst0__I2;
  wire [0:0] Mux10x1_inst0__I3;
  wire [0:0] Mux10x1_inst0__I4;
  wire [0:0] Mux10x1_inst0__I5;
  wire [0:0] Mux10x1_inst0__I6;
  wire [0:0] Mux10x1_inst0__I7;
  wire [0:0] Mux10x1_inst0__I8;
  wire [0:0] Mux10x1_inst0__I9;
  wire [0:0] Mux10x1_inst0__O;
  wire [3:0] Mux10x1_inst0__S;
  Mux10x1 Mux10x1_inst0(
    .I0(Mux10x1_inst0__I0),
    .I1(Mux10x1_inst0__I1),
    .I2(Mux10x1_inst0__I2),
    .I3(Mux10x1_inst0__I3),
    .I4(Mux10x1_inst0__I4),
    .I5(Mux10x1_inst0__I5),
    .I6(Mux10x1_inst0__I6),
    .I7(Mux10x1_inst0__I7),
    .I8(Mux10x1_inst0__I8),
    .I9(Mux10x1_inst0__I9),
    .O(Mux10x1_inst0__O),
    .S(Mux10x1_inst0__S)
  );

  assign Mux10x1_inst0__I0[0:0] = I_0[0:0];

  assign Mux10x1_inst0__I1[0:0] = I_1[0:0];

  assign Mux10x1_inst0__I2[0:0] = I_2[0:0];

  assign Mux10x1_inst0__I3[0:0] = I_3[0:0];

  assign Mux10x1_inst0__I4[0:0] = I_4[0:0];

  assign Mux10x1_inst0__I5[0:0] = I_5[0:0];

  assign Mux10x1_inst0__I6[0:0] = I_6[0:0];

  assign Mux10x1_inst0__I7[0:0] = I_7[0:0];

  assign Mux10x1_inst0__I8[0:0] = I_8[0:0];

  assign Mux10x1_inst0__I9[0:0] = I_9[0:0];

  assign O[0:0] = Mux10x1_inst0__O[0:0];

  assign Mux10x1_inst0__S[3:0] = S[3:0];


endmodule  // MuxWrapper_10_1

module Decode68 (
  input [7:0] I,
  output  O
);


  // Instancing generated Module: coreir.const(width:8)
  wire [7:0] const_6_8__out;
  coreir_const #(.value(8'h06),.width(8)) const_6_8(
    .out(const_6_8__out)
  );

  // Instancing generated Module: coreir.eq(width:8)
  wire [7:0] coreir_eq_8_inst0__in0;
  wire [7:0] coreir_eq_8_inst0__in1;
  wire  coreir_eq_8_inst0__out;
  coreir_eq #(.width(8)) coreir_eq_8_inst0(
    .in0(coreir_eq_8_inst0__in0),
    .in1(coreir_eq_8_inst0__in1),
    .out(coreir_eq_8_inst0__out)
  );

  assign coreir_eq_8_inst0__in1[7:0] = const_6_8__out[7:0];

  assign coreir_eq_8_inst0__in0[7:0] = I[7:0];

  assign O = coreir_eq_8_inst0__out;


endmodule  // Decode68

module Decode58 (
  input [7:0] I,
  output  O
);


  // Instancing generated Module: coreir.const(width:8)
  wire [7:0] const_5_8__out;
  coreir_const #(.value(8'h05),.width(8)) const_5_8(
    .out(const_5_8__out)
  );

  // Instancing generated Module: coreir.eq(width:8)
  wire [7:0] coreir_eq_8_inst0__in0;
  wire [7:0] coreir_eq_8_inst0__in1;
  wire  coreir_eq_8_inst0__out;
  coreir_eq #(.width(8)) coreir_eq_8_inst0(
    .in0(coreir_eq_8_inst0__in0),
    .in1(coreir_eq_8_inst0__in1),
    .out(coreir_eq_8_inst0__out)
  );

  assign coreir_eq_8_inst0__in1[7:0] = const_5_8__out[7:0];

  assign coreir_eq_8_inst0__in0[7:0] = I[7:0];

  assign O = coreir_eq_8_inst0__out;


endmodule  // Decode58

module Decode48 (
  input [7:0] I,
  output  O
);


  // Instancing generated Module: coreir.const(width:8)
  wire [7:0] const_4_8__out;
  coreir_const #(.value(8'h04),.width(8)) const_4_8(
    .out(const_4_8__out)
  );

  // Instancing generated Module: coreir.eq(width:8)
  wire [7:0] coreir_eq_8_inst0__in0;
  wire [7:0] coreir_eq_8_inst0__in1;
  wire  coreir_eq_8_inst0__out;
  coreir_eq #(.width(8)) coreir_eq_8_inst0(
    .in0(coreir_eq_8_inst0__in0),
    .in1(coreir_eq_8_inst0__in1),
    .out(coreir_eq_8_inst0__out)
  );

  assign coreir_eq_8_inst0__in1[7:0] = const_4_8__out[7:0];

  assign coreir_eq_8_inst0__in0[7:0] = I[7:0];

  assign O = coreir_eq_8_inst0__out;


endmodule  // Decode48

module Decode38 (
  input [7:0] I,
  output  O
);


  // Instancing generated Module: coreir.const(width:8)
  wire [7:0] const_3_8__out;
  coreir_const #(.value(8'h03),.width(8)) const_3_8(
    .out(const_3_8__out)
  );

  // Instancing generated Module: coreir.eq(width:8)
  wire [7:0] coreir_eq_8_inst0__in0;
  wire [7:0] coreir_eq_8_inst0__in1;
  wire  coreir_eq_8_inst0__out;
  coreir_eq #(.width(8)) coreir_eq_8_inst0(
    .in0(coreir_eq_8_inst0__in0),
    .in1(coreir_eq_8_inst0__in1),
    .out(coreir_eq_8_inst0__out)
  );

  assign coreir_eq_8_inst0__in1[7:0] = const_3_8__out[7:0];

  assign coreir_eq_8_inst0__in0[7:0] = I[7:0];

  assign O = coreir_eq_8_inst0__out;


endmodule  // Decode38

module Decode28 (
  input [7:0] I,
  output  O
);


  // Instancing generated Module: coreir.const(width:8)
  wire [7:0] const_2_8__out;
  coreir_const #(.value(8'h02),.width(8)) const_2_8(
    .out(const_2_8__out)
  );

  // Instancing generated Module: coreir.eq(width:8)
  wire [7:0] coreir_eq_8_inst0__in0;
  wire [7:0] coreir_eq_8_inst0__in1;
  wire  coreir_eq_8_inst0__out;
  coreir_eq #(.width(8)) coreir_eq_8_inst0(
    .in0(coreir_eq_8_inst0__in0),
    .in1(coreir_eq_8_inst0__in1),
    .out(coreir_eq_8_inst0__out)
  );

  assign coreir_eq_8_inst0__in1[7:0] = const_2_8__out[7:0];

  assign coreir_eq_8_inst0__in0[7:0] = I[7:0];

  assign O = coreir_eq_8_inst0__out;


endmodule  // Decode28

module Decode18 (
  input [7:0] I,
  output  O
);


  // Instancing generated Module: coreir.const(width:8)
  wire [7:0] const_1_8__out;
  coreir_const #(.value(8'h01),.width(8)) const_1_8(
    .out(const_1_8__out)
  );

  // Instancing generated Module: coreir.eq(width:8)
  wire [7:0] coreir_eq_8_inst0__in0;
  wire [7:0] coreir_eq_8_inst0__in1;
  wire  coreir_eq_8_inst0__out;
  coreir_eq #(.width(8)) coreir_eq_8_inst0(
    .in0(coreir_eq_8_inst0__in0),
    .in1(coreir_eq_8_inst0__in1),
    .out(coreir_eq_8_inst0__out)
  );

  assign coreir_eq_8_inst0__in1[7:0] = const_1_8__out[7:0];

  assign coreir_eq_8_inst0__in0[7:0] = I[7:0];

  assign O = coreir_eq_8_inst0__out;


endmodule  // Decode18

module Decode08 (
  input [7:0] I,
  output  O
);


  // Instancing generated Module: coreir.const(width:8)
  wire [7:0] const_0_8__out;
  coreir_const #(.value(8'h00),.width(8)) const_0_8(
    .out(const_0_8__out)
  );

  // Instancing generated Module: coreir.eq(width:8)
  wire [7:0] coreir_eq_8_inst0__in0;
  wire [7:0] coreir_eq_8_inst0__in1;
  wire  coreir_eq_8_inst0__out;
  coreir_eq #(.width(8)) coreir_eq_8_inst0(
    .in0(coreir_eq_8_inst0__in0),
    .in1(coreir_eq_8_inst0__in1),
    .out(coreir_eq_8_inst0__out)
  );

  assign coreir_eq_8_inst0__in1[7:0] = const_0_8__out[7:0];

  assign coreir_eq_8_inst0__in0[7:0] = I[7:0];

  assign O = coreir_eq_8_inst0__out;


endmodule  // Decode08

module ConfigRegister_4_8_32_0 (
  output [3:0] O,
  input  clk,
  input [7:0] config_addr,
  input [31:0] config_data,
  input  config_en,
  input  reset
);


  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_4_inst0__ASYNCRESET;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_4_inst0__CE;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_4_inst0__CLK;
  wire [3:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_4_inst0__I;
  wire [3:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_4_inst0__O;
  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_4 Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_4_inst0(
    .ASYNCRESET(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_4_inst0__ASYNCRESET),
    .CE(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_4_inst0__CE),
    .CLK(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_4_inst0__CLK),
    .I(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_4_inst0__I),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_4_inst0__O)
  );

  wire  and_inst0__in0;
  wire  and_inst0__in1;
  wire  and_inst0__out;
  corebit_and and_inst0(
    .in0(and_inst0__in0),
    .in1(and_inst0__in1),
    .out(and_inst0__out)
  );

  // Instancing generated Module: coreir.const(width:8)
  wire [7:0] const_0_8__out;
  coreir_const #(.value(8'h00),.width(8)) const_0_8(
    .out(const_0_8__out)
  );

  // Instancing generated Module: coreir.eq(width:8)
  wire [7:0] coreir_eq_8_inst0__in0;
  wire [7:0] coreir_eq_8_inst0__in1;
  wire  coreir_eq_8_inst0__out;
  coreir_eq #(.width(8)) coreir_eq_8_inst0(
    .in0(coreir_eq_8_inst0__in0),
    .in1(coreir_eq_8_inst0__in1),
    .out(coreir_eq_8_inst0__out)
  );

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_4_inst0__ASYNCRESET = reset;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_4_inst0__CE = and_inst0__out;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_4_inst0__CLK = clk;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_4_inst0__I[0] = config_data[0];

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_4_inst0__I[1] = config_data[1];

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_4_inst0__I[2] = config_data[2];

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_4_inst0__I[3] = config_data[3];

  assign O[3:0] = Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_4_inst0__O[3:0];

  assign and_inst0__in0 = coreir_eq_8_inst0__out;

  assign and_inst0__in1 = config_en;

  assign coreir_eq_8_inst0__in1[7:0] = const_0_8__out[7:0];

  assign coreir_eq_8_inst0__in0[7:0] = config_addr[7:0];


endmodule  // ConfigRegister_4_8_32_0

module ConfigRegister_2_8_32_8 (
  output [1:0] O,
  input  clk,
  input [7:0] config_addr,
  input [31:0] config_data,
  input  config_en,
  input  reset
);


  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK;
  wire [1:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I;
  wire [1:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O;
  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2 Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0(
    .ASYNCRESET(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET),
    .CE(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE),
    .CLK(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK),
    .I(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O)
  );

  wire  and_inst0__in0;
  wire  and_inst0__in1;
  wire  and_inst0__out;
  corebit_and and_inst0(
    .in0(and_inst0__in0),
    .in1(and_inst0__in1),
    .out(and_inst0__out)
  );

  // Instancing generated Module: coreir.const(width:8)
  wire [7:0] const_8_8__out;
  coreir_const #(.value(8'h08),.width(8)) const_8_8(
    .out(const_8_8__out)
  );

  // Instancing generated Module: coreir.eq(width:8)
  wire [7:0] coreir_eq_8_inst0__in0;
  wire [7:0] coreir_eq_8_inst0__in1;
  wire  coreir_eq_8_inst0__out;
  coreir_eq #(.width(8)) coreir_eq_8_inst0(
    .in0(coreir_eq_8_inst0__in0),
    .in1(coreir_eq_8_inst0__in1),
    .out(coreir_eq_8_inst0__out)
  );

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET = reset;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE = and_inst0__out;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK = clk;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I[0] = config_data[0];

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I[1] = config_data[1];

  assign O[1:0] = Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O[1:0];

  assign and_inst0__in0 = coreir_eq_8_inst0__out;

  assign and_inst0__in1 = config_en;

  assign coreir_eq_8_inst0__in1[7:0] = const_8_8__out[7:0];

  assign coreir_eq_8_inst0__in0[7:0] = config_addr[7:0];


endmodule  // ConfigRegister_2_8_32_8

module ConfigRegister_2_8_32_78 (
  output [1:0] O,
  input  clk,
  input [7:0] config_addr,
  input [31:0] config_data,
  input  config_en,
  input  reset
);


  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK;
  wire [1:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I;
  wire [1:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O;
  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2 Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0(
    .ASYNCRESET(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET),
    .CE(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE),
    .CLK(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK),
    .I(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O)
  );

  wire  and_inst0__in0;
  wire  and_inst0__in1;
  wire  and_inst0__out;
  corebit_and and_inst0(
    .in0(and_inst0__in0),
    .in1(and_inst0__in1),
    .out(and_inst0__out)
  );

  // Instancing generated Module: coreir.const(width:8)
  wire [7:0] const_78_8__out;
  coreir_const #(.value(8'h4e),.width(8)) const_78_8(
    .out(const_78_8__out)
  );

  // Instancing generated Module: coreir.eq(width:8)
  wire [7:0] coreir_eq_8_inst0__in0;
  wire [7:0] coreir_eq_8_inst0__in1;
  wire  coreir_eq_8_inst0__out;
  coreir_eq #(.width(8)) coreir_eq_8_inst0(
    .in0(coreir_eq_8_inst0__in0),
    .in1(coreir_eq_8_inst0__in1),
    .out(coreir_eq_8_inst0__out)
  );

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET = reset;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE = and_inst0__out;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK = clk;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I[0] = config_data[0];

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I[1] = config_data[1];

  assign O[1:0] = Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O[1:0];

  assign and_inst0__in0 = coreir_eq_8_inst0__out;

  assign and_inst0__in1 = config_en;

  assign coreir_eq_8_inst0__in1[7:0] = const_78_8__out[7:0];

  assign coreir_eq_8_inst0__in0[7:0] = config_addr[7:0];


endmodule  // ConfigRegister_2_8_32_78

module ConfigRegister_2_8_32_76 (
  output [1:0] O,
  input  clk,
  input [7:0] config_addr,
  input [31:0] config_data,
  input  config_en,
  input  reset
);


  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK;
  wire [1:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I;
  wire [1:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O;
  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2 Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0(
    .ASYNCRESET(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET),
    .CE(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE),
    .CLK(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK),
    .I(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O)
  );

  wire  and_inst0__in0;
  wire  and_inst0__in1;
  wire  and_inst0__out;
  corebit_and and_inst0(
    .in0(and_inst0__in0),
    .in1(and_inst0__in1),
    .out(and_inst0__out)
  );

  // Instancing generated Module: coreir.const(width:8)
  wire [7:0] const_76_8__out;
  coreir_const #(.value(8'h4c),.width(8)) const_76_8(
    .out(const_76_8__out)
  );

  // Instancing generated Module: coreir.eq(width:8)
  wire [7:0] coreir_eq_8_inst0__in0;
  wire [7:0] coreir_eq_8_inst0__in1;
  wire  coreir_eq_8_inst0__out;
  coreir_eq #(.width(8)) coreir_eq_8_inst0(
    .in0(coreir_eq_8_inst0__in0),
    .in1(coreir_eq_8_inst0__in1),
    .out(coreir_eq_8_inst0__out)
  );

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET = reset;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE = and_inst0__out;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK = clk;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I[0] = config_data[0];

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I[1] = config_data[1];

  assign O[1:0] = Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O[1:0];

  assign and_inst0__in0 = coreir_eq_8_inst0__out;

  assign and_inst0__in1 = config_en;

  assign coreir_eq_8_inst0__in1[7:0] = const_76_8__out[7:0];

  assign coreir_eq_8_inst0__in0[7:0] = config_addr[7:0];


endmodule  // ConfigRegister_2_8_32_76

module ConfigRegister_2_8_32_74 (
  output [1:0] O,
  input  clk,
  input [7:0] config_addr,
  input [31:0] config_data,
  input  config_en,
  input  reset
);


  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK;
  wire [1:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I;
  wire [1:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O;
  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2 Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0(
    .ASYNCRESET(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET),
    .CE(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE),
    .CLK(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK),
    .I(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O)
  );

  wire  and_inst0__in0;
  wire  and_inst0__in1;
  wire  and_inst0__out;
  corebit_and and_inst0(
    .in0(and_inst0__in0),
    .in1(and_inst0__in1),
    .out(and_inst0__out)
  );

  // Instancing generated Module: coreir.const(width:8)
  wire [7:0] const_74_8__out;
  coreir_const #(.value(8'h4a),.width(8)) const_74_8(
    .out(const_74_8__out)
  );

  // Instancing generated Module: coreir.eq(width:8)
  wire [7:0] coreir_eq_8_inst0__in0;
  wire [7:0] coreir_eq_8_inst0__in1;
  wire  coreir_eq_8_inst0__out;
  coreir_eq #(.width(8)) coreir_eq_8_inst0(
    .in0(coreir_eq_8_inst0__in0),
    .in1(coreir_eq_8_inst0__in1),
    .out(coreir_eq_8_inst0__out)
  );

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET = reset;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE = and_inst0__out;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK = clk;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I[0] = config_data[0];

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I[1] = config_data[1];

  assign O[1:0] = Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O[1:0];

  assign and_inst0__in0 = coreir_eq_8_inst0__out;

  assign and_inst0__in1 = config_en;

  assign coreir_eq_8_inst0__in1[7:0] = const_74_8__out[7:0];

  assign coreir_eq_8_inst0__in0[7:0] = config_addr[7:0];


endmodule  // ConfigRegister_2_8_32_74

module ConfigRegister_2_8_32_72 (
  output [1:0] O,
  input  clk,
  input [7:0] config_addr,
  input [31:0] config_data,
  input  config_en,
  input  reset
);


  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK;
  wire [1:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I;
  wire [1:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O;
  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2 Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0(
    .ASYNCRESET(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET),
    .CE(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE),
    .CLK(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK),
    .I(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O)
  );

  wire  and_inst0__in0;
  wire  and_inst0__in1;
  wire  and_inst0__out;
  corebit_and and_inst0(
    .in0(and_inst0__in0),
    .in1(and_inst0__in1),
    .out(and_inst0__out)
  );

  // Instancing generated Module: coreir.const(width:8)
  wire [7:0] const_72_8__out;
  coreir_const #(.value(8'h48),.width(8)) const_72_8(
    .out(const_72_8__out)
  );

  // Instancing generated Module: coreir.eq(width:8)
  wire [7:0] coreir_eq_8_inst0__in0;
  wire [7:0] coreir_eq_8_inst0__in1;
  wire  coreir_eq_8_inst0__out;
  coreir_eq #(.width(8)) coreir_eq_8_inst0(
    .in0(coreir_eq_8_inst0__in0),
    .in1(coreir_eq_8_inst0__in1),
    .out(coreir_eq_8_inst0__out)
  );

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET = reset;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE = and_inst0__out;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK = clk;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I[0] = config_data[0];

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I[1] = config_data[1];

  assign O[1:0] = Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O[1:0];

  assign and_inst0__in0 = coreir_eq_8_inst0__out;

  assign and_inst0__in1 = config_en;

  assign coreir_eq_8_inst0__in1[7:0] = const_72_8__out[7:0];

  assign coreir_eq_8_inst0__in0[7:0] = config_addr[7:0];


endmodule  // ConfigRegister_2_8_32_72

module ConfigRegister_2_8_32_70 (
  output [1:0] O,
  input  clk,
  input [7:0] config_addr,
  input [31:0] config_data,
  input  config_en,
  input  reset
);


  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK;
  wire [1:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I;
  wire [1:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O;
  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2 Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0(
    .ASYNCRESET(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET),
    .CE(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE),
    .CLK(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK),
    .I(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O)
  );

  wire  and_inst0__in0;
  wire  and_inst0__in1;
  wire  and_inst0__out;
  corebit_and and_inst0(
    .in0(and_inst0__in0),
    .in1(and_inst0__in1),
    .out(and_inst0__out)
  );

  // Instancing generated Module: coreir.const(width:8)
  wire [7:0] const_70_8__out;
  coreir_const #(.value(8'h46),.width(8)) const_70_8(
    .out(const_70_8__out)
  );

  // Instancing generated Module: coreir.eq(width:8)
  wire [7:0] coreir_eq_8_inst0__in0;
  wire [7:0] coreir_eq_8_inst0__in1;
  wire  coreir_eq_8_inst0__out;
  coreir_eq #(.width(8)) coreir_eq_8_inst0(
    .in0(coreir_eq_8_inst0__in0),
    .in1(coreir_eq_8_inst0__in1),
    .out(coreir_eq_8_inst0__out)
  );

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET = reset;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE = and_inst0__out;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK = clk;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I[0] = config_data[0];

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I[1] = config_data[1];

  assign O[1:0] = Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O[1:0];

  assign and_inst0__in0 = coreir_eq_8_inst0__out;

  assign and_inst0__in1 = config_en;

  assign coreir_eq_8_inst0__in1[7:0] = const_70_8__out[7:0];

  assign coreir_eq_8_inst0__in0[7:0] = config_addr[7:0];


endmodule  // ConfigRegister_2_8_32_70

module ConfigRegister_2_8_32_68 (
  output [1:0] O,
  input  clk,
  input [7:0] config_addr,
  input [31:0] config_data,
  input  config_en,
  input  reset
);


  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK;
  wire [1:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I;
  wire [1:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O;
  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2 Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0(
    .ASYNCRESET(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET),
    .CE(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE),
    .CLK(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK),
    .I(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O)
  );

  wire  and_inst0__in0;
  wire  and_inst0__in1;
  wire  and_inst0__out;
  corebit_and and_inst0(
    .in0(and_inst0__in0),
    .in1(and_inst0__in1),
    .out(and_inst0__out)
  );

  // Instancing generated Module: coreir.const(width:8)
  wire [7:0] const_68_8__out;
  coreir_const #(.value(8'h44),.width(8)) const_68_8(
    .out(const_68_8__out)
  );

  // Instancing generated Module: coreir.eq(width:8)
  wire [7:0] coreir_eq_8_inst0__in0;
  wire [7:0] coreir_eq_8_inst0__in1;
  wire  coreir_eq_8_inst0__out;
  coreir_eq #(.width(8)) coreir_eq_8_inst0(
    .in0(coreir_eq_8_inst0__in0),
    .in1(coreir_eq_8_inst0__in1),
    .out(coreir_eq_8_inst0__out)
  );

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET = reset;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE = and_inst0__out;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK = clk;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I[0] = config_data[0];

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I[1] = config_data[1];

  assign O[1:0] = Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O[1:0];

  assign and_inst0__in0 = coreir_eq_8_inst0__out;

  assign and_inst0__in1 = config_en;

  assign coreir_eq_8_inst0__in1[7:0] = const_68_8__out[7:0];

  assign coreir_eq_8_inst0__in0[7:0] = config_addr[7:0];


endmodule  // ConfigRegister_2_8_32_68

module ConfigRegister_2_8_32_66 (
  output [1:0] O,
  input  clk,
  input [7:0] config_addr,
  input [31:0] config_data,
  input  config_en,
  input  reset
);


  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK;
  wire [1:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I;
  wire [1:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O;
  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2 Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0(
    .ASYNCRESET(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET),
    .CE(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE),
    .CLK(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK),
    .I(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O)
  );

  wire  and_inst0__in0;
  wire  and_inst0__in1;
  wire  and_inst0__out;
  corebit_and and_inst0(
    .in0(and_inst0__in0),
    .in1(and_inst0__in1),
    .out(and_inst0__out)
  );

  // Instancing generated Module: coreir.const(width:8)
  wire [7:0] const_66_8__out;
  coreir_const #(.value(8'h42),.width(8)) const_66_8(
    .out(const_66_8__out)
  );

  // Instancing generated Module: coreir.eq(width:8)
  wire [7:0] coreir_eq_8_inst0__in0;
  wire [7:0] coreir_eq_8_inst0__in1;
  wire  coreir_eq_8_inst0__out;
  coreir_eq #(.width(8)) coreir_eq_8_inst0(
    .in0(coreir_eq_8_inst0__in0),
    .in1(coreir_eq_8_inst0__in1),
    .out(coreir_eq_8_inst0__out)
  );

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET = reset;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE = and_inst0__out;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK = clk;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I[0] = config_data[0];

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I[1] = config_data[1];

  assign O[1:0] = Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O[1:0];

  assign and_inst0__in0 = coreir_eq_8_inst0__out;

  assign and_inst0__in1 = config_en;

  assign coreir_eq_8_inst0__in1[7:0] = const_66_8__out[7:0];

  assign coreir_eq_8_inst0__in0[7:0] = config_addr[7:0];


endmodule  // ConfigRegister_2_8_32_66

module ConfigRegister_2_8_32_64 (
  output [1:0] O,
  input  clk,
  input [7:0] config_addr,
  input [31:0] config_data,
  input  config_en,
  input  reset
);


  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK;
  wire [1:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I;
  wire [1:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O;
  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2 Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0(
    .ASYNCRESET(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET),
    .CE(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE),
    .CLK(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK),
    .I(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O)
  );

  wire  and_inst0__in0;
  wire  and_inst0__in1;
  wire  and_inst0__out;
  corebit_and and_inst0(
    .in0(and_inst0__in0),
    .in1(and_inst0__in1),
    .out(and_inst0__out)
  );

  // Instancing generated Module: coreir.const(width:8)
  wire [7:0] const_64_8__out;
  coreir_const #(.value(8'h40),.width(8)) const_64_8(
    .out(const_64_8__out)
  );

  // Instancing generated Module: coreir.eq(width:8)
  wire [7:0] coreir_eq_8_inst0__in0;
  wire [7:0] coreir_eq_8_inst0__in1;
  wire  coreir_eq_8_inst0__out;
  coreir_eq #(.width(8)) coreir_eq_8_inst0(
    .in0(coreir_eq_8_inst0__in0),
    .in1(coreir_eq_8_inst0__in1),
    .out(coreir_eq_8_inst0__out)
  );

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET = reset;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE = and_inst0__out;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK = clk;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I[0] = config_data[0];

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I[1] = config_data[1];

  assign O[1:0] = Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O[1:0];

  assign and_inst0__in0 = coreir_eq_8_inst0__out;

  assign and_inst0__in1 = config_en;

  assign coreir_eq_8_inst0__in1[7:0] = const_64_8__out[7:0];

  assign coreir_eq_8_inst0__in0[7:0] = config_addr[7:0];


endmodule  // ConfigRegister_2_8_32_64

module ConfigRegister_2_8_32_62 (
  output [1:0] O,
  input  clk,
  input [7:0] config_addr,
  input [31:0] config_data,
  input  config_en,
  input  reset
);


  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK;
  wire [1:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I;
  wire [1:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O;
  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2 Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0(
    .ASYNCRESET(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET),
    .CE(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE),
    .CLK(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK),
    .I(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O)
  );

  wire  and_inst0__in0;
  wire  and_inst0__in1;
  wire  and_inst0__out;
  corebit_and and_inst0(
    .in0(and_inst0__in0),
    .in1(and_inst0__in1),
    .out(and_inst0__out)
  );

  // Instancing generated Module: coreir.const(width:8)
  wire [7:0] const_62_8__out;
  coreir_const #(.value(8'h3e),.width(8)) const_62_8(
    .out(const_62_8__out)
  );

  // Instancing generated Module: coreir.eq(width:8)
  wire [7:0] coreir_eq_8_inst0__in0;
  wire [7:0] coreir_eq_8_inst0__in1;
  wire  coreir_eq_8_inst0__out;
  coreir_eq #(.width(8)) coreir_eq_8_inst0(
    .in0(coreir_eq_8_inst0__in0),
    .in1(coreir_eq_8_inst0__in1),
    .out(coreir_eq_8_inst0__out)
  );

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET = reset;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE = and_inst0__out;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK = clk;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I[0] = config_data[0];

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I[1] = config_data[1];

  assign O[1:0] = Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O[1:0];

  assign and_inst0__in0 = coreir_eq_8_inst0__out;

  assign and_inst0__in1 = config_en;

  assign coreir_eq_8_inst0__in1[7:0] = const_62_8__out[7:0];

  assign coreir_eq_8_inst0__in0[7:0] = config_addr[7:0];


endmodule  // ConfigRegister_2_8_32_62

module ConfigRegister_2_8_32_60 (
  output [1:0] O,
  input  clk,
  input [7:0] config_addr,
  input [31:0] config_data,
  input  config_en,
  input  reset
);


  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK;
  wire [1:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I;
  wire [1:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O;
  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2 Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0(
    .ASYNCRESET(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET),
    .CE(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE),
    .CLK(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK),
    .I(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O)
  );

  wire  and_inst0__in0;
  wire  and_inst0__in1;
  wire  and_inst0__out;
  corebit_and and_inst0(
    .in0(and_inst0__in0),
    .in1(and_inst0__in1),
    .out(and_inst0__out)
  );

  // Instancing generated Module: coreir.const(width:8)
  wire [7:0] const_60_8__out;
  coreir_const #(.value(8'h3c),.width(8)) const_60_8(
    .out(const_60_8__out)
  );

  // Instancing generated Module: coreir.eq(width:8)
  wire [7:0] coreir_eq_8_inst0__in0;
  wire [7:0] coreir_eq_8_inst0__in1;
  wire  coreir_eq_8_inst0__out;
  coreir_eq #(.width(8)) coreir_eq_8_inst0(
    .in0(coreir_eq_8_inst0__in0),
    .in1(coreir_eq_8_inst0__in1),
    .out(coreir_eq_8_inst0__out)
  );

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET = reset;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE = and_inst0__out;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK = clk;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I[0] = config_data[0];

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I[1] = config_data[1];

  assign O[1:0] = Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O[1:0];

  assign and_inst0__in0 = coreir_eq_8_inst0__out;

  assign and_inst0__in1 = config_en;

  assign coreir_eq_8_inst0__in1[7:0] = const_60_8__out[7:0];

  assign coreir_eq_8_inst0__in0[7:0] = config_addr[7:0];


endmodule  // ConfigRegister_2_8_32_60

module ConfigRegister_2_8_32_6 (
  output [1:0] O,
  input  clk,
  input [7:0] config_addr,
  input [31:0] config_data,
  input  config_en,
  input  reset
);


  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK;
  wire [1:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I;
  wire [1:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O;
  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2 Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0(
    .ASYNCRESET(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET),
    .CE(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE),
    .CLK(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK),
    .I(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O)
  );

  wire  and_inst0__in0;
  wire  and_inst0__in1;
  wire  and_inst0__out;
  corebit_and and_inst0(
    .in0(and_inst0__in0),
    .in1(and_inst0__in1),
    .out(and_inst0__out)
  );

  // Instancing generated Module: coreir.const(width:8)
  wire [7:0] const_6_8__out;
  coreir_const #(.value(8'h06),.width(8)) const_6_8(
    .out(const_6_8__out)
  );

  // Instancing generated Module: coreir.eq(width:8)
  wire [7:0] coreir_eq_8_inst0__in0;
  wire [7:0] coreir_eq_8_inst0__in1;
  wire  coreir_eq_8_inst0__out;
  coreir_eq #(.width(8)) coreir_eq_8_inst0(
    .in0(coreir_eq_8_inst0__in0),
    .in1(coreir_eq_8_inst0__in1),
    .out(coreir_eq_8_inst0__out)
  );

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET = reset;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE = and_inst0__out;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK = clk;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I[0] = config_data[0];

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I[1] = config_data[1];

  assign O[1:0] = Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O[1:0];

  assign and_inst0__in0 = coreir_eq_8_inst0__out;

  assign and_inst0__in1 = config_en;

  assign coreir_eq_8_inst0__in1[7:0] = const_6_8__out[7:0];

  assign coreir_eq_8_inst0__in0[7:0] = config_addr[7:0];


endmodule  // ConfigRegister_2_8_32_6

module ConfigRegister_2_8_32_58 (
  output [1:0] O,
  input  clk,
  input [7:0] config_addr,
  input [31:0] config_data,
  input  config_en,
  input  reset
);


  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK;
  wire [1:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I;
  wire [1:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O;
  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2 Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0(
    .ASYNCRESET(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET),
    .CE(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE),
    .CLK(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK),
    .I(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O)
  );

  wire  and_inst0__in0;
  wire  and_inst0__in1;
  wire  and_inst0__out;
  corebit_and and_inst0(
    .in0(and_inst0__in0),
    .in1(and_inst0__in1),
    .out(and_inst0__out)
  );

  // Instancing generated Module: coreir.const(width:8)
  wire [7:0] const_58_8__out;
  coreir_const #(.value(8'h3a),.width(8)) const_58_8(
    .out(const_58_8__out)
  );

  // Instancing generated Module: coreir.eq(width:8)
  wire [7:0] coreir_eq_8_inst0__in0;
  wire [7:0] coreir_eq_8_inst0__in1;
  wire  coreir_eq_8_inst0__out;
  coreir_eq #(.width(8)) coreir_eq_8_inst0(
    .in0(coreir_eq_8_inst0__in0),
    .in1(coreir_eq_8_inst0__in1),
    .out(coreir_eq_8_inst0__out)
  );

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET = reset;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE = and_inst0__out;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK = clk;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I[0] = config_data[0];

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I[1] = config_data[1];

  assign O[1:0] = Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O[1:0];

  assign and_inst0__in0 = coreir_eq_8_inst0__out;

  assign and_inst0__in1 = config_en;

  assign coreir_eq_8_inst0__in1[7:0] = const_58_8__out[7:0];

  assign coreir_eq_8_inst0__in0[7:0] = config_addr[7:0];


endmodule  // ConfigRegister_2_8_32_58

module ConfigRegister_2_8_32_56 (
  output [1:0] O,
  input  clk,
  input [7:0] config_addr,
  input [31:0] config_data,
  input  config_en,
  input  reset
);


  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK;
  wire [1:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I;
  wire [1:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O;
  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2 Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0(
    .ASYNCRESET(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET),
    .CE(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE),
    .CLK(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK),
    .I(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O)
  );

  wire  and_inst0__in0;
  wire  and_inst0__in1;
  wire  and_inst0__out;
  corebit_and and_inst0(
    .in0(and_inst0__in0),
    .in1(and_inst0__in1),
    .out(and_inst0__out)
  );

  // Instancing generated Module: coreir.const(width:8)
  wire [7:0] const_56_8__out;
  coreir_const #(.value(8'h38),.width(8)) const_56_8(
    .out(const_56_8__out)
  );

  // Instancing generated Module: coreir.eq(width:8)
  wire [7:0] coreir_eq_8_inst0__in0;
  wire [7:0] coreir_eq_8_inst0__in1;
  wire  coreir_eq_8_inst0__out;
  coreir_eq #(.width(8)) coreir_eq_8_inst0(
    .in0(coreir_eq_8_inst0__in0),
    .in1(coreir_eq_8_inst0__in1),
    .out(coreir_eq_8_inst0__out)
  );

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET = reset;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE = and_inst0__out;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK = clk;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I[0] = config_data[0];

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I[1] = config_data[1];

  assign O[1:0] = Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O[1:0];

  assign and_inst0__in0 = coreir_eq_8_inst0__out;

  assign and_inst0__in1 = config_en;

  assign coreir_eq_8_inst0__in1[7:0] = const_56_8__out[7:0];

  assign coreir_eq_8_inst0__in0[7:0] = config_addr[7:0];


endmodule  // ConfigRegister_2_8_32_56

module ConfigRegister_2_8_32_54 (
  output [1:0] O,
  input  clk,
  input [7:0] config_addr,
  input [31:0] config_data,
  input  config_en,
  input  reset
);


  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK;
  wire [1:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I;
  wire [1:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O;
  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2 Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0(
    .ASYNCRESET(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET),
    .CE(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE),
    .CLK(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK),
    .I(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O)
  );

  wire  and_inst0__in0;
  wire  and_inst0__in1;
  wire  and_inst0__out;
  corebit_and and_inst0(
    .in0(and_inst0__in0),
    .in1(and_inst0__in1),
    .out(and_inst0__out)
  );

  // Instancing generated Module: coreir.const(width:8)
  wire [7:0] const_54_8__out;
  coreir_const #(.value(8'h36),.width(8)) const_54_8(
    .out(const_54_8__out)
  );

  // Instancing generated Module: coreir.eq(width:8)
  wire [7:0] coreir_eq_8_inst0__in0;
  wire [7:0] coreir_eq_8_inst0__in1;
  wire  coreir_eq_8_inst0__out;
  coreir_eq #(.width(8)) coreir_eq_8_inst0(
    .in0(coreir_eq_8_inst0__in0),
    .in1(coreir_eq_8_inst0__in1),
    .out(coreir_eq_8_inst0__out)
  );

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET = reset;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE = and_inst0__out;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK = clk;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I[0] = config_data[0];

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I[1] = config_data[1];

  assign O[1:0] = Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O[1:0];

  assign and_inst0__in0 = coreir_eq_8_inst0__out;

  assign and_inst0__in1 = config_en;

  assign coreir_eq_8_inst0__in1[7:0] = const_54_8__out[7:0];

  assign coreir_eq_8_inst0__in0[7:0] = config_addr[7:0];


endmodule  // ConfigRegister_2_8_32_54

module ConfigRegister_2_8_32_52 (
  output [1:0] O,
  input  clk,
  input [7:0] config_addr,
  input [31:0] config_data,
  input  config_en,
  input  reset
);


  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK;
  wire [1:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I;
  wire [1:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O;
  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2 Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0(
    .ASYNCRESET(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET),
    .CE(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE),
    .CLK(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK),
    .I(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O)
  );

  wire  and_inst0__in0;
  wire  and_inst0__in1;
  wire  and_inst0__out;
  corebit_and and_inst0(
    .in0(and_inst0__in0),
    .in1(and_inst0__in1),
    .out(and_inst0__out)
  );

  // Instancing generated Module: coreir.const(width:8)
  wire [7:0] const_52_8__out;
  coreir_const #(.value(8'h34),.width(8)) const_52_8(
    .out(const_52_8__out)
  );

  // Instancing generated Module: coreir.eq(width:8)
  wire [7:0] coreir_eq_8_inst0__in0;
  wire [7:0] coreir_eq_8_inst0__in1;
  wire  coreir_eq_8_inst0__out;
  coreir_eq #(.width(8)) coreir_eq_8_inst0(
    .in0(coreir_eq_8_inst0__in0),
    .in1(coreir_eq_8_inst0__in1),
    .out(coreir_eq_8_inst0__out)
  );

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET = reset;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE = and_inst0__out;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK = clk;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I[0] = config_data[0];

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I[1] = config_data[1];

  assign O[1:0] = Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O[1:0];

  assign and_inst0__in0 = coreir_eq_8_inst0__out;

  assign and_inst0__in1 = config_en;

  assign coreir_eq_8_inst0__in1[7:0] = const_52_8__out[7:0];

  assign coreir_eq_8_inst0__in0[7:0] = config_addr[7:0];


endmodule  // ConfigRegister_2_8_32_52

module ConfigRegister_2_8_32_50 (
  output [1:0] O,
  input  clk,
  input [7:0] config_addr,
  input [31:0] config_data,
  input  config_en,
  input  reset
);


  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK;
  wire [1:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I;
  wire [1:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O;
  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2 Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0(
    .ASYNCRESET(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET),
    .CE(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE),
    .CLK(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK),
    .I(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O)
  );

  wire  and_inst0__in0;
  wire  and_inst0__in1;
  wire  and_inst0__out;
  corebit_and and_inst0(
    .in0(and_inst0__in0),
    .in1(and_inst0__in1),
    .out(and_inst0__out)
  );

  // Instancing generated Module: coreir.const(width:8)
  wire [7:0] const_50_8__out;
  coreir_const #(.value(8'h32),.width(8)) const_50_8(
    .out(const_50_8__out)
  );

  // Instancing generated Module: coreir.eq(width:8)
  wire [7:0] coreir_eq_8_inst0__in0;
  wire [7:0] coreir_eq_8_inst0__in1;
  wire  coreir_eq_8_inst0__out;
  coreir_eq #(.width(8)) coreir_eq_8_inst0(
    .in0(coreir_eq_8_inst0__in0),
    .in1(coreir_eq_8_inst0__in1),
    .out(coreir_eq_8_inst0__out)
  );

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET = reset;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE = and_inst0__out;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK = clk;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I[0] = config_data[0];

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I[1] = config_data[1];

  assign O[1:0] = Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O[1:0];

  assign and_inst0__in0 = coreir_eq_8_inst0__out;

  assign and_inst0__in1 = config_en;

  assign coreir_eq_8_inst0__in1[7:0] = const_50_8__out[7:0];

  assign coreir_eq_8_inst0__in0[7:0] = config_addr[7:0];


endmodule  // ConfigRegister_2_8_32_50

module ConfigRegister_2_8_32_48 (
  output [1:0] O,
  input  clk,
  input [7:0] config_addr,
  input [31:0] config_data,
  input  config_en,
  input  reset
);


  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK;
  wire [1:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I;
  wire [1:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O;
  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2 Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0(
    .ASYNCRESET(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET),
    .CE(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE),
    .CLK(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK),
    .I(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O)
  );

  wire  and_inst0__in0;
  wire  and_inst0__in1;
  wire  and_inst0__out;
  corebit_and and_inst0(
    .in0(and_inst0__in0),
    .in1(and_inst0__in1),
    .out(and_inst0__out)
  );

  // Instancing generated Module: coreir.const(width:8)
  wire [7:0] const_48_8__out;
  coreir_const #(.value(8'h30),.width(8)) const_48_8(
    .out(const_48_8__out)
  );

  // Instancing generated Module: coreir.eq(width:8)
  wire [7:0] coreir_eq_8_inst0__in0;
  wire [7:0] coreir_eq_8_inst0__in1;
  wire  coreir_eq_8_inst0__out;
  coreir_eq #(.width(8)) coreir_eq_8_inst0(
    .in0(coreir_eq_8_inst0__in0),
    .in1(coreir_eq_8_inst0__in1),
    .out(coreir_eq_8_inst0__out)
  );

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET = reset;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE = and_inst0__out;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK = clk;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I[0] = config_data[0];

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I[1] = config_data[1];

  assign O[1:0] = Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O[1:0];

  assign and_inst0__in0 = coreir_eq_8_inst0__out;

  assign and_inst0__in1 = config_en;

  assign coreir_eq_8_inst0__in1[7:0] = const_48_8__out[7:0];

  assign coreir_eq_8_inst0__in0[7:0] = config_addr[7:0];


endmodule  // ConfigRegister_2_8_32_48

module ConfigRegister_2_8_32_46 (
  output [1:0] O,
  input  clk,
  input [7:0] config_addr,
  input [31:0] config_data,
  input  config_en,
  input  reset
);


  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK;
  wire [1:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I;
  wire [1:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O;
  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2 Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0(
    .ASYNCRESET(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET),
    .CE(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE),
    .CLK(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK),
    .I(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O)
  );

  wire  and_inst0__in0;
  wire  and_inst0__in1;
  wire  and_inst0__out;
  corebit_and and_inst0(
    .in0(and_inst0__in0),
    .in1(and_inst0__in1),
    .out(and_inst0__out)
  );

  // Instancing generated Module: coreir.const(width:8)
  wire [7:0] const_46_8__out;
  coreir_const #(.value(8'h2e),.width(8)) const_46_8(
    .out(const_46_8__out)
  );

  // Instancing generated Module: coreir.eq(width:8)
  wire [7:0] coreir_eq_8_inst0__in0;
  wire [7:0] coreir_eq_8_inst0__in1;
  wire  coreir_eq_8_inst0__out;
  coreir_eq #(.width(8)) coreir_eq_8_inst0(
    .in0(coreir_eq_8_inst0__in0),
    .in1(coreir_eq_8_inst0__in1),
    .out(coreir_eq_8_inst0__out)
  );

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET = reset;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE = and_inst0__out;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK = clk;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I[0] = config_data[0];

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I[1] = config_data[1];

  assign O[1:0] = Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O[1:0];

  assign and_inst0__in0 = coreir_eq_8_inst0__out;

  assign and_inst0__in1 = config_en;

  assign coreir_eq_8_inst0__in1[7:0] = const_46_8__out[7:0];

  assign coreir_eq_8_inst0__in0[7:0] = config_addr[7:0];


endmodule  // ConfigRegister_2_8_32_46

module ConfigRegister_2_8_32_44 (
  output [1:0] O,
  input  clk,
  input [7:0] config_addr,
  input [31:0] config_data,
  input  config_en,
  input  reset
);


  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK;
  wire [1:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I;
  wire [1:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O;
  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2 Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0(
    .ASYNCRESET(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET),
    .CE(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE),
    .CLK(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK),
    .I(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O)
  );

  wire  and_inst0__in0;
  wire  and_inst0__in1;
  wire  and_inst0__out;
  corebit_and and_inst0(
    .in0(and_inst0__in0),
    .in1(and_inst0__in1),
    .out(and_inst0__out)
  );

  // Instancing generated Module: coreir.const(width:8)
  wire [7:0] const_44_8__out;
  coreir_const #(.value(8'h2c),.width(8)) const_44_8(
    .out(const_44_8__out)
  );

  // Instancing generated Module: coreir.eq(width:8)
  wire [7:0] coreir_eq_8_inst0__in0;
  wire [7:0] coreir_eq_8_inst0__in1;
  wire  coreir_eq_8_inst0__out;
  coreir_eq #(.width(8)) coreir_eq_8_inst0(
    .in0(coreir_eq_8_inst0__in0),
    .in1(coreir_eq_8_inst0__in1),
    .out(coreir_eq_8_inst0__out)
  );

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET = reset;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE = and_inst0__out;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK = clk;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I[0] = config_data[0];

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I[1] = config_data[1];

  assign O[1:0] = Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O[1:0];

  assign and_inst0__in0 = coreir_eq_8_inst0__out;

  assign and_inst0__in1 = config_en;

  assign coreir_eq_8_inst0__in1[7:0] = const_44_8__out[7:0];

  assign coreir_eq_8_inst0__in0[7:0] = config_addr[7:0];


endmodule  // ConfigRegister_2_8_32_44

module ConfigRegister_2_8_32_42 (
  output [1:0] O,
  input  clk,
  input [7:0] config_addr,
  input [31:0] config_data,
  input  config_en,
  input  reset
);


  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK;
  wire [1:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I;
  wire [1:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O;
  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2 Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0(
    .ASYNCRESET(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET),
    .CE(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE),
    .CLK(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK),
    .I(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O)
  );

  wire  and_inst0__in0;
  wire  and_inst0__in1;
  wire  and_inst0__out;
  corebit_and and_inst0(
    .in0(and_inst0__in0),
    .in1(and_inst0__in1),
    .out(and_inst0__out)
  );

  // Instancing generated Module: coreir.const(width:8)
  wire [7:0] const_42_8__out;
  coreir_const #(.value(8'h2a),.width(8)) const_42_8(
    .out(const_42_8__out)
  );

  // Instancing generated Module: coreir.eq(width:8)
  wire [7:0] coreir_eq_8_inst0__in0;
  wire [7:0] coreir_eq_8_inst0__in1;
  wire  coreir_eq_8_inst0__out;
  coreir_eq #(.width(8)) coreir_eq_8_inst0(
    .in0(coreir_eq_8_inst0__in0),
    .in1(coreir_eq_8_inst0__in1),
    .out(coreir_eq_8_inst0__out)
  );

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET = reset;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE = and_inst0__out;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK = clk;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I[0] = config_data[0];

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I[1] = config_data[1];

  assign O[1:0] = Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O[1:0];

  assign and_inst0__in0 = coreir_eq_8_inst0__out;

  assign and_inst0__in1 = config_en;

  assign coreir_eq_8_inst0__in1[7:0] = const_42_8__out[7:0];

  assign coreir_eq_8_inst0__in0[7:0] = config_addr[7:0];


endmodule  // ConfigRegister_2_8_32_42

module ConfigRegister_2_8_32_40 (
  output [1:0] O,
  input  clk,
  input [7:0] config_addr,
  input [31:0] config_data,
  input  config_en,
  input  reset
);


  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK;
  wire [1:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I;
  wire [1:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O;
  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2 Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0(
    .ASYNCRESET(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET),
    .CE(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE),
    .CLK(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK),
    .I(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O)
  );

  wire  and_inst0__in0;
  wire  and_inst0__in1;
  wire  and_inst0__out;
  corebit_and and_inst0(
    .in0(and_inst0__in0),
    .in1(and_inst0__in1),
    .out(and_inst0__out)
  );

  // Instancing generated Module: coreir.const(width:8)
  wire [7:0] const_40_8__out;
  coreir_const #(.value(8'h28),.width(8)) const_40_8(
    .out(const_40_8__out)
  );

  // Instancing generated Module: coreir.eq(width:8)
  wire [7:0] coreir_eq_8_inst0__in0;
  wire [7:0] coreir_eq_8_inst0__in1;
  wire  coreir_eq_8_inst0__out;
  coreir_eq #(.width(8)) coreir_eq_8_inst0(
    .in0(coreir_eq_8_inst0__in0),
    .in1(coreir_eq_8_inst0__in1),
    .out(coreir_eq_8_inst0__out)
  );

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET = reset;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE = and_inst0__out;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK = clk;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I[0] = config_data[0];

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I[1] = config_data[1];

  assign O[1:0] = Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O[1:0];

  assign and_inst0__in0 = coreir_eq_8_inst0__out;

  assign and_inst0__in1 = config_en;

  assign coreir_eq_8_inst0__in1[7:0] = const_40_8__out[7:0];

  assign coreir_eq_8_inst0__in0[7:0] = config_addr[7:0];


endmodule  // ConfigRegister_2_8_32_40

module ConfigRegister_2_8_32_4 (
  output [1:0] O,
  input  clk,
  input [7:0] config_addr,
  input [31:0] config_data,
  input  config_en,
  input  reset
);


  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK;
  wire [1:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I;
  wire [1:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O;
  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2 Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0(
    .ASYNCRESET(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET),
    .CE(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE),
    .CLK(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK),
    .I(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O)
  );

  wire  and_inst0__in0;
  wire  and_inst0__in1;
  wire  and_inst0__out;
  corebit_and and_inst0(
    .in0(and_inst0__in0),
    .in1(and_inst0__in1),
    .out(and_inst0__out)
  );

  // Instancing generated Module: coreir.const(width:8)
  wire [7:0] const_4_8__out;
  coreir_const #(.value(8'h04),.width(8)) const_4_8(
    .out(const_4_8__out)
  );

  // Instancing generated Module: coreir.eq(width:8)
  wire [7:0] coreir_eq_8_inst0__in0;
  wire [7:0] coreir_eq_8_inst0__in1;
  wire  coreir_eq_8_inst0__out;
  coreir_eq #(.width(8)) coreir_eq_8_inst0(
    .in0(coreir_eq_8_inst0__in0),
    .in1(coreir_eq_8_inst0__in1),
    .out(coreir_eq_8_inst0__out)
  );

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET = reset;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE = and_inst0__out;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK = clk;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I[0] = config_data[0];

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I[1] = config_data[1];

  assign O[1:0] = Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O[1:0];

  assign and_inst0__in0 = coreir_eq_8_inst0__out;

  assign and_inst0__in1 = config_en;

  assign coreir_eq_8_inst0__in1[7:0] = const_4_8__out[7:0];

  assign coreir_eq_8_inst0__in0[7:0] = config_addr[7:0];


endmodule  // ConfigRegister_2_8_32_4

module ConfigRegister_2_8_32_38 (
  output [1:0] O,
  input  clk,
  input [7:0] config_addr,
  input [31:0] config_data,
  input  config_en,
  input  reset
);


  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK;
  wire [1:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I;
  wire [1:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O;
  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2 Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0(
    .ASYNCRESET(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET),
    .CE(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE),
    .CLK(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK),
    .I(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O)
  );

  wire  and_inst0__in0;
  wire  and_inst0__in1;
  wire  and_inst0__out;
  corebit_and and_inst0(
    .in0(and_inst0__in0),
    .in1(and_inst0__in1),
    .out(and_inst0__out)
  );

  // Instancing generated Module: coreir.const(width:8)
  wire [7:0] const_38_8__out;
  coreir_const #(.value(8'h26),.width(8)) const_38_8(
    .out(const_38_8__out)
  );

  // Instancing generated Module: coreir.eq(width:8)
  wire [7:0] coreir_eq_8_inst0__in0;
  wire [7:0] coreir_eq_8_inst0__in1;
  wire  coreir_eq_8_inst0__out;
  coreir_eq #(.width(8)) coreir_eq_8_inst0(
    .in0(coreir_eq_8_inst0__in0),
    .in1(coreir_eq_8_inst0__in1),
    .out(coreir_eq_8_inst0__out)
  );

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET = reset;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE = and_inst0__out;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK = clk;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I[0] = config_data[0];

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I[1] = config_data[1];

  assign O[1:0] = Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O[1:0];

  assign and_inst0__in0 = coreir_eq_8_inst0__out;

  assign and_inst0__in1 = config_en;

  assign coreir_eq_8_inst0__in1[7:0] = const_38_8__out[7:0];

  assign coreir_eq_8_inst0__in0[7:0] = config_addr[7:0];


endmodule  // ConfigRegister_2_8_32_38

module ConfigRegister_2_8_32_36 (
  output [1:0] O,
  input  clk,
  input [7:0] config_addr,
  input [31:0] config_data,
  input  config_en,
  input  reset
);


  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK;
  wire [1:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I;
  wire [1:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O;
  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2 Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0(
    .ASYNCRESET(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET),
    .CE(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE),
    .CLK(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK),
    .I(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O)
  );

  wire  and_inst0__in0;
  wire  and_inst0__in1;
  wire  and_inst0__out;
  corebit_and and_inst0(
    .in0(and_inst0__in0),
    .in1(and_inst0__in1),
    .out(and_inst0__out)
  );

  // Instancing generated Module: coreir.const(width:8)
  wire [7:0] const_36_8__out;
  coreir_const #(.value(8'h24),.width(8)) const_36_8(
    .out(const_36_8__out)
  );

  // Instancing generated Module: coreir.eq(width:8)
  wire [7:0] coreir_eq_8_inst0__in0;
  wire [7:0] coreir_eq_8_inst0__in1;
  wire  coreir_eq_8_inst0__out;
  coreir_eq #(.width(8)) coreir_eq_8_inst0(
    .in0(coreir_eq_8_inst0__in0),
    .in1(coreir_eq_8_inst0__in1),
    .out(coreir_eq_8_inst0__out)
  );

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET = reset;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE = and_inst0__out;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK = clk;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I[0] = config_data[0];

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I[1] = config_data[1];

  assign O[1:0] = Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O[1:0];

  assign and_inst0__in0 = coreir_eq_8_inst0__out;

  assign and_inst0__in1 = config_en;

  assign coreir_eq_8_inst0__in1[7:0] = const_36_8__out[7:0];

  assign coreir_eq_8_inst0__in0[7:0] = config_addr[7:0];


endmodule  // ConfigRegister_2_8_32_36

module ConfigRegister_2_8_32_34 (
  output [1:0] O,
  input  clk,
  input [7:0] config_addr,
  input [31:0] config_data,
  input  config_en,
  input  reset
);


  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK;
  wire [1:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I;
  wire [1:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O;
  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2 Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0(
    .ASYNCRESET(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET),
    .CE(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE),
    .CLK(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK),
    .I(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O)
  );

  wire  and_inst0__in0;
  wire  and_inst0__in1;
  wire  and_inst0__out;
  corebit_and and_inst0(
    .in0(and_inst0__in0),
    .in1(and_inst0__in1),
    .out(and_inst0__out)
  );

  // Instancing generated Module: coreir.const(width:8)
  wire [7:0] const_34_8__out;
  coreir_const #(.value(8'h22),.width(8)) const_34_8(
    .out(const_34_8__out)
  );

  // Instancing generated Module: coreir.eq(width:8)
  wire [7:0] coreir_eq_8_inst0__in0;
  wire [7:0] coreir_eq_8_inst0__in1;
  wire  coreir_eq_8_inst0__out;
  coreir_eq #(.width(8)) coreir_eq_8_inst0(
    .in0(coreir_eq_8_inst0__in0),
    .in1(coreir_eq_8_inst0__in1),
    .out(coreir_eq_8_inst0__out)
  );

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET = reset;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE = and_inst0__out;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK = clk;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I[0] = config_data[0];

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I[1] = config_data[1];

  assign O[1:0] = Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O[1:0];

  assign and_inst0__in0 = coreir_eq_8_inst0__out;

  assign and_inst0__in1 = config_en;

  assign coreir_eq_8_inst0__in1[7:0] = const_34_8__out[7:0];

  assign coreir_eq_8_inst0__in0[7:0] = config_addr[7:0];


endmodule  // ConfigRegister_2_8_32_34

module ConfigRegister_2_8_32_32 (
  output [1:0] O,
  input  clk,
  input [7:0] config_addr,
  input [31:0] config_data,
  input  config_en,
  input  reset
);


  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK;
  wire [1:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I;
  wire [1:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O;
  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2 Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0(
    .ASYNCRESET(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET),
    .CE(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE),
    .CLK(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK),
    .I(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O)
  );

  wire  and_inst0__in0;
  wire  and_inst0__in1;
  wire  and_inst0__out;
  corebit_and and_inst0(
    .in0(and_inst0__in0),
    .in1(and_inst0__in1),
    .out(and_inst0__out)
  );

  // Instancing generated Module: coreir.const(width:8)
  wire [7:0] const_32_8__out;
  coreir_const #(.value(8'h20),.width(8)) const_32_8(
    .out(const_32_8__out)
  );

  // Instancing generated Module: coreir.eq(width:8)
  wire [7:0] coreir_eq_8_inst0__in0;
  wire [7:0] coreir_eq_8_inst0__in1;
  wire  coreir_eq_8_inst0__out;
  coreir_eq #(.width(8)) coreir_eq_8_inst0(
    .in0(coreir_eq_8_inst0__in0),
    .in1(coreir_eq_8_inst0__in1),
    .out(coreir_eq_8_inst0__out)
  );

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET = reset;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE = and_inst0__out;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK = clk;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I[0] = config_data[0];

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I[1] = config_data[1];

  assign O[1:0] = Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O[1:0];

  assign and_inst0__in0 = coreir_eq_8_inst0__out;

  assign and_inst0__in1 = config_en;

  assign coreir_eq_8_inst0__in1[7:0] = const_32_8__out[7:0];

  assign coreir_eq_8_inst0__in0[7:0] = config_addr[7:0];


endmodule  // ConfigRegister_2_8_32_32

module ConfigRegister_2_8_32_30 (
  output [1:0] O,
  input  clk,
  input [7:0] config_addr,
  input [31:0] config_data,
  input  config_en,
  input  reset
);


  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK;
  wire [1:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I;
  wire [1:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O;
  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2 Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0(
    .ASYNCRESET(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET),
    .CE(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE),
    .CLK(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK),
    .I(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O)
  );

  wire  and_inst0__in0;
  wire  and_inst0__in1;
  wire  and_inst0__out;
  corebit_and and_inst0(
    .in0(and_inst0__in0),
    .in1(and_inst0__in1),
    .out(and_inst0__out)
  );

  // Instancing generated Module: coreir.const(width:8)
  wire [7:0] const_30_8__out;
  coreir_const #(.value(8'h1e),.width(8)) const_30_8(
    .out(const_30_8__out)
  );

  // Instancing generated Module: coreir.eq(width:8)
  wire [7:0] coreir_eq_8_inst0__in0;
  wire [7:0] coreir_eq_8_inst0__in1;
  wire  coreir_eq_8_inst0__out;
  coreir_eq #(.width(8)) coreir_eq_8_inst0(
    .in0(coreir_eq_8_inst0__in0),
    .in1(coreir_eq_8_inst0__in1),
    .out(coreir_eq_8_inst0__out)
  );

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET = reset;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE = and_inst0__out;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK = clk;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I[0] = config_data[0];

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I[1] = config_data[1];

  assign O[1:0] = Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O[1:0];

  assign and_inst0__in0 = coreir_eq_8_inst0__out;

  assign and_inst0__in1 = config_en;

  assign coreir_eq_8_inst0__in1[7:0] = const_30_8__out[7:0];

  assign coreir_eq_8_inst0__in0[7:0] = config_addr[7:0];


endmodule  // ConfigRegister_2_8_32_30

module ConfigRegister_2_8_32_28 (
  output [1:0] O,
  input  clk,
  input [7:0] config_addr,
  input [31:0] config_data,
  input  config_en,
  input  reset
);


  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK;
  wire [1:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I;
  wire [1:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O;
  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2 Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0(
    .ASYNCRESET(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET),
    .CE(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE),
    .CLK(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK),
    .I(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O)
  );

  wire  and_inst0__in0;
  wire  and_inst0__in1;
  wire  and_inst0__out;
  corebit_and and_inst0(
    .in0(and_inst0__in0),
    .in1(and_inst0__in1),
    .out(and_inst0__out)
  );

  // Instancing generated Module: coreir.const(width:8)
  wire [7:0] const_28_8__out;
  coreir_const #(.value(8'h1c),.width(8)) const_28_8(
    .out(const_28_8__out)
  );

  // Instancing generated Module: coreir.eq(width:8)
  wire [7:0] coreir_eq_8_inst0__in0;
  wire [7:0] coreir_eq_8_inst0__in1;
  wire  coreir_eq_8_inst0__out;
  coreir_eq #(.width(8)) coreir_eq_8_inst0(
    .in0(coreir_eq_8_inst0__in0),
    .in1(coreir_eq_8_inst0__in1),
    .out(coreir_eq_8_inst0__out)
  );

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET = reset;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE = and_inst0__out;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK = clk;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I[0] = config_data[0];

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I[1] = config_data[1];

  assign O[1:0] = Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O[1:0];

  assign and_inst0__in0 = coreir_eq_8_inst0__out;

  assign and_inst0__in1 = config_en;

  assign coreir_eq_8_inst0__in1[7:0] = const_28_8__out[7:0];

  assign coreir_eq_8_inst0__in0[7:0] = config_addr[7:0];


endmodule  // ConfigRegister_2_8_32_28

module ConfigRegister_2_8_32_26 (
  output [1:0] O,
  input  clk,
  input [7:0] config_addr,
  input [31:0] config_data,
  input  config_en,
  input  reset
);


  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK;
  wire [1:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I;
  wire [1:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O;
  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2 Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0(
    .ASYNCRESET(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET),
    .CE(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE),
    .CLK(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK),
    .I(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O)
  );

  wire  and_inst0__in0;
  wire  and_inst0__in1;
  wire  and_inst0__out;
  corebit_and and_inst0(
    .in0(and_inst0__in0),
    .in1(and_inst0__in1),
    .out(and_inst0__out)
  );

  // Instancing generated Module: coreir.const(width:8)
  wire [7:0] const_26_8__out;
  coreir_const #(.value(8'h1a),.width(8)) const_26_8(
    .out(const_26_8__out)
  );

  // Instancing generated Module: coreir.eq(width:8)
  wire [7:0] coreir_eq_8_inst0__in0;
  wire [7:0] coreir_eq_8_inst0__in1;
  wire  coreir_eq_8_inst0__out;
  coreir_eq #(.width(8)) coreir_eq_8_inst0(
    .in0(coreir_eq_8_inst0__in0),
    .in1(coreir_eq_8_inst0__in1),
    .out(coreir_eq_8_inst0__out)
  );

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET = reset;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE = and_inst0__out;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK = clk;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I[0] = config_data[0];

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I[1] = config_data[1];

  assign O[1:0] = Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O[1:0];

  assign and_inst0__in0 = coreir_eq_8_inst0__out;

  assign and_inst0__in1 = config_en;

  assign coreir_eq_8_inst0__in1[7:0] = const_26_8__out[7:0];

  assign coreir_eq_8_inst0__in0[7:0] = config_addr[7:0];


endmodule  // ConfigRegister_2_8_32_26

module ConfigRegister_2_8_32_24 (
  output [1:0] O,
  input  clk,
  input [7:0] config_addr,
  input [31:0] config_data,
  input  config_en,
  input  reset
);


  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK;
  wire [1:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I;
  wire [1:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O;
  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2 Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0(
    .ASYNCRESET(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET),
    .CE(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE),
    .CLK(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK),
    .I(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O)
  );

  wire  and_inst0__in0;
  wire  and_inst0__in1;
  wire  and_inst0__out;
  corebit_and and_inst0(
    .in0(and_inst0__in0),
    .in1(and_inst0__in1),
    .out(and_inst0__out)
  );

  // Instancing generated Module: coreir.const(width:8)
  wire [7:0] const_24_8__out;
  coreir_const #(.value(8'h18),.width(8)) const_24_8(
    .out(const_24_8__out)
  );

  // Instancing generated Module: coreir.eq(width:8)
  wire [7:0] coreir_eq_8_inst0__in0;
  wire [7:0] coreir_eq_8_inst0__in1;
  wire  coreir_eq_8_inst0__out;
  coreir_eq #(.width(8)) coreir_eq_8_inst0(
    .in0(coreir_eq_8_inst0__in0),
    .in1(coreir_eq_8_inst0__in1),
    .out(coreir_eq_8_inst0__out)
  );

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET = reset;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE = and_inst0__out;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK = clk;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I[0] = config_data[0];

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I[1] = config_data[1];

  assign O[1:0] = Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O[1:0];

  assign and_inst0__in0 = coreir_eq_8_inst0__out;

  assign and_inst0__in1 = config_en;

  assign coreir_eq_8_inst0__in1[7:0] = const_24_8__out[7:0];

  assign coreir_eq_8_inst0__in0[7:0] = config_addr[7:0];


endmodule  // ConfigRegister_2_8_32_24

module ConfigRegister_2_8_32_22 (
  output [1:0] O,
  input  clk,
  input [7:0] config_addr,
  input [31:0] config_data,
  input  config_en,
  input  reset
);


  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK;
  wire [1:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I;
  wire [1:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O;
  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2 Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0(
    .ASYNCRESET(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET),
    .CE(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE),
    .CLK(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK),
    .I(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O)
  );

  wire  and_inst0__in0;
  wire  and_inst0__in1;
  wire  and_inst0__out;
  corebit_and and_inst0(
    .in0(and_inst0__in0),
    .in1(and_inst0__in1),
    .out(and_inst0__out)
  );

  // Instancing generated Module: coreir.const(width:8)
  wire [7:0] const_22_8__out;
  coreir_const #(.value(8'h16),.width(8)) const_22_8(
    .out(const_22_8__out)
  );

  // Instancing generated Module: coreir.eq(width:8)
  wire [7:0] coreir_eq_8_inst0__in0;
  wire [7:0] coreir_eq_8_inst0__in1;
  wire  coreir_eq_8_inst0__out;
  coreir_eq #(.width(8)) coreir_eq_8_inst0(
    .in0(coreir_eq_8_inst0__in0),
    .in1(coreir_eq_8_inst0__in1),
    .out(coreir_eq_8_inst0__out)
  );

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET = reset;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE = and_inst0__out;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK = clk;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I[0] = config_data[0];

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I[1] = config_data[1];

  assign O[1:0] = Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O[1:0];

  assign and_inst0__in0 = coreir_eq_8_inst0__out;

  assign and_inst0__in1 = config_en;

  assign coreir_eq_8_inst0__in1[7:0] = const_22_8__out[7:0];

  assign coreir_eq_8_inst0__in0[7:0] = config_addr[7:0];


endmodule  // ConfigRegister_2_8_32_22

module ConfigRegister_2_8_32_20 (
  output [1:0] O,
  input  clk,
  input [7:0] config_addr,
  input [31:0] config_data,
  input  config_en,
  input  reset
);


  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK;
  wire [1:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I;
  wire [1:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O;
  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2 Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0(
    .ASYNCRESET(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET),
    .CE(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE),
    .CLK(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK),
    .I(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O)
  );

  wire  and_inst0__in0;
  wire  and_inst0__in1;
  wire  and_inst0__out;
  corebit_and and_inst0(
    .in0(and_inst0__in0),
    .in1(and_inst0__in1),
    .out(and_inst0__out)
  );

  // Instancing generated Module: coreir.const(width:8)
  wire [7:0] const_20_8__out;
  coreir_const #(.value(8'h14),.width(8)) const_20_8(
    .out(const_20_8__out)
  );

  // Instancing generated Module: coreir.eq(width:8)
  wire [7:0] coreir_eq_8_inst0__in0;
  wire [7:0] coreir_eq_8_inst0__in1;
  wire  coreir_eq_8_inst0__out;
  coreir_eq #(.width(8)) coreir_eq_8_inst0(
    .in0(coreir_eq_8_inst0__in0),
    .in1(coreir_eq_8_inst0__in1),
    .out(coreir_eq_8_inst0__out)
  );

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET = reset;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE = and_inst0__out;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK = clk;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I[0] = config_data[0];

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I[1] = config_data[1];

  assign O[1:0] = Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O[1:0];

  assign and_inst0__in0 = coreir_eq_8_inst0__out;

  assign and_inst0__in1 = config_en;

  assign coreir_eq_8_inst0__in1[7:0] = const_20_8__out[7:0];

  assign coreir_eq_8_inst0__in0[7:0] = config_addr[7:0];


endmodule  // ConfigRegister_2_8_32_20

module ConfigRegister_2_8_32_2 (
  output [1:0] O,
  input  clk,
  input [7:0] config_addr,
  input [31:0] config_data,
  input  config_en,
  input  reset
);


  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK;
  wire [1:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I;
  wire [1:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O;
  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2 Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0(
    .ASYNCRESET(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET),
    .CE(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE),
    .CLK(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK),
    .I(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O)
  );

  wire  and_inst0__in0;
  wire  and_inst0__in1;
  wire  and_inst0__out;
  corebit_and and_inst0(
    .in0(and_inst0__in0),
    .in1(and_inst0__in1),
    .out(and_inst0__out)
  );

  // Instancing generated Module: coreir.const(width:8)
  wire [7:0] const_2_8__out;
  coreir_const #(.value(8'h02),.width(8)) const_2_8(
    .out(const_2_8__out)
  );

  // Instancing generated Module: coreir.eq(width:8)
  wire [7:0] coreir_eq_8_inst0__in0;
  wire [7:0] coreir_eq_8_inst0__in1;
  wire  coreir_eq_8_inst0__out;
  coreir_eq #(.width(8)) coreir_eq_8_inst0(
    .in0(coreir_eq_8_inst0__in0),
    .in1(coreir_eq_8_inst0__in1),
    .out(coreir_eq_8_inst0__out)
  );

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET = reset;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE = and_inst0__out;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK = clk;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I[0] = config_data[0];

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I[1] = config_data[1];

  assign O[1:0] = Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O[1:0];

  assign and_inst0__in0 = coreir_eq_8_inst0__out;

  assign and_inst0__in1 = config_en;

  assign coreir_eq_8_inst0__in1[7:0] = const_2_8__out[7:0];

  assign coreir_eq_8_inst0__in0[7:0] = config_addr[7:0];


endmodule  // ConfigRegister_2_8_32_2

module ConfigRegister_2_8_32_18 (
  output [1:0] O,
  input  clk,
  input [7:0] config_addr,
  input [31:0] config_data,
  input  config_en,
  input  reset
);


  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK;
  wire [1:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I;
  wire [1:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O;
  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2 Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0(
    .ASYNCRESET(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET),
    .CE(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE),
    .CLK(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK),
    .I(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O)
  );

  wire  and_inst0__in0;
  wire  and_inst0__in1;
  wire  and_inst0__out;
  corebit_and and_inst0(
    .in0(and_inst0__in0),
    .in1(and_inst0__in1),
    .out(and_inst0__out)
  );

  // Instancing generated Module: coreir.const(width:8)
  wire [7:0] const_18_8__out;
  coreir_const #(.value(8'h12),.width(8)) const_18_8(
    .out(const_18_8__out)
  );

  // Instancing generated Module: coreir.eq(width:8)
  wire [7:0] coreir_eq_8_inst0__in0;
  wire [7:0] coreir_eq_8_inst0__in1;
  wire  coreir_eq_8_inst0__out;
  coreir_eq #(.width(8)) coreir_eq_8_inst0(
    .in0(coreir_eq_8_inst0__in0),
    .in1(coreir_eq_8_inst0__in1),
    .out(coreir_eq_8_inst0__out)
  );

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET = reset;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE = and_inst0__out;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK = clk;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I[0] = config_data[0];

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I[1] = config_data[1];

  assign O[1:0] = Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O[1:0];

  assign and_inst0__in0 = coreir_eq_8_inst0__out;

  assign and_inst0__in1 = config_en;

  assign coreir_eq_8_inst0__in1[7:0] = const_18_8__out[7:0];

  assign coreir_eq_8_inst0__in0[7:0] = config_addr[7:0];


endmodule  // ConfigRegister_2_8_32_18

module ConfigRegister_2_8_32_16 (
  output [1:0] O,
  input  clk,
  input [7:0] config_addr,
  input [31:0] config_data,
  input  config_en,
  input  reset
);


  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK;
  wire [1:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I;
  wire [1:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O;
  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2 Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0(
    .ASYNCRESET(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET),
    .CE(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE),
    .CLK(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK),
    .I(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O)
  );

  wire  and_inst0__in0;
  wire  and_inst0__in1;
  wire  and_inst0__out;
  corebit_and and_inst0(
    .in0(and_inst0__in0),
    .in1(and_inst0__in1),
    .out(and_inst0__out)
  );

  // Instancing generated Module: coreir.const(width:8)
  wire [7:0] const_16_8__out;
  coreir_const #(.value(8'h10),.width(8)) const_16_8(
    .out(const_16_8__out)
  );

  // Instancing generated Module: coreir.eq(width:8)
  wire [7:0] coreir_eq_8_inst0__in0;
  wire [7:0] coreir_eq_8_inst0__in1;
  wire  coreir_eq_8_inst0__out;
  coreir_eq #(.width(8)) coreir_eq_8_inst0(
    .in0(coreir_eq_8_inst0__in0),
    .in1(coreir_eq_8_inst0__in1),
    .out(coreir_eq_8_inst0__out)
  );

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET = reset;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE = and_inst0__out;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK = clk;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I[0] = config_data[0];

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I[1] = config_data[1];

  assign O[1:0] = Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O[1:0];

  assign and_inst0__in0 = coreir_eq_8_inst0__out;

  assign and_inst0__in1 = config_en;

  assign coreir_eq_8_inst0__in1[7:0] = const_16_8__out[7:0];

  assign coreir_eq_8_inst0__in0[7:0] = config_addr[7:0];


endmodule  // ConfigRegister_2_8_32_16

module ConfigRegister_2_8_32_14 (
  output [1:0] O,
  input  clk,
  input [7:0] config_addr,
  input [31:0] config_data,
  input  config_en,
  input  reset
);


  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK;
  wire [1:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I;
  wire [1:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O;
  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2 Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0(
    .ASYNCRESET(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET),
    .CE(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE),
    .CLK(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK),
    .I(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O)
  );

  wire  and_inst0__in0;
  wire  and_inst0__in1;
  wire  and_inst0__out;
  corebit_and and_inst0(
    .in0(and_inst0__in0),
    .in1(and_inst0__in1),
    .out(and_inst0__out)
  );

  // Instancing generated Module: coreir.const(width:8)
  wire [7:0] const_14_8__out;
  coreir_const #(.value(8'h0e),.width(8)) const_14_8(
    .out(const_14_8__out)
  );

  // Instancing generated Module: coreir.eq(width:8)
  wire [7:0] coreir_eq_8_inst0__in0;
  wire [7:0] coreir_eq_8_inst0__in1;
  wire  coreir_eq_8_inst0__out;
  coreir_eq #(.width(8)) coreir_eq_8_inst0(
    .in0(coreir_eq_8_inst0__in0),
    .in1(coreir_eq_8_inst0__in1),
    .out(coreir_eq_8_inst0__out)
  );

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET = reset;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE = and_inst0__out;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK = clk;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I[0] = config_data[0];

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I[1] = config_data[1];

  assign O[1:0] = Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O[1:0];

  assign and_inst0__in0 = coreir_eq_8_inst0__out;

  assign and_inst0__in1 = config_en;

  assign coreir_eq_8_inst0__in1[7:0] = const_14_8__out[7:0];

  assign coreir_eq_8_inst0__in0[7:0] = config_addr[7:0];


endmodule  // ConfigRegister_2_8_32_14

module ConfigRegister_2_8_32_12 (
  output [1:0] O,
  input  clk,
  input [7:0] config_addr,
  input [31:0] config_data,
  input  config_en,
  input  reset
);


  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK;
  wire [1:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I;
  wire [1:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O;
  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2 Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0(
    .ASYNCRESET(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET),
    .CE(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE),
    .CLK(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK),
    .I(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O)
  );

  wire  and_inst0__in0;
  wire  and_inst0__in1;
  wire  and_inst0__out;
  corebit_and and_inst0(
    .in0(and_inst0__in0),
    .in1(and_inst0__in1),
    .out(and_inst0__out)
  );

  // Instancing generated Module: coreir.const(width:8)
  wire [7:0] const_12_8__out;
  coreir_const #(.value(8'h0c),.width(8)) const_12_8(
    .out(const_12_8__out)
  );

  // Instancing generated Module: coreir.eq(width:8)
  wire [7:0] coreir_eq_8_inst0__in0;
  wire [7:0] coreir_eq_8_inst0__in1;
  wire  coreir_eq_8_inst0__out;
  coreir_eq #(.width(8)) coreir_eq_8_inst0(
    .in0(coreir_eq_8_inst0__in0),
    .in1(coreir_eq_8_inst0__in1),
    .out(coreir_eq_8_inst0__out)
  );

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET = reset;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE = and_inst0__out;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK = clk;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I[0] = config_data[0];

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I[1] = config_data[1];

  assign O[1:0] = Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O[1:0];

  assign and_inst0__in0 = coreir_eq_8_inst0__out;

  assign and_inst0__in1 = config_en;

  assign coreir_eq_8_inst0__in1[7:0] = const_12_8__out[7:0];

  assign coreir_eq_8_inst0__in0[7:0] = config_addr[7:0];


endmodule  // ConfigRegister_2_8_32_12

module ConfigRegister_2_8_32_10 (
  output [1:0] O,
  input  clk,
  input [7:0] config_addr,
  input [31:0] config_data,
  input  config_en,
  input  reset
);


  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK;
  wire [1:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I;
  wire [1:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O;
  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2 Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0(
    .ASYNCRESET(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET),
    .CE(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE),
    .CLK(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK),
    .I(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O)
  );

  wire  and_inst0__in0;
  wire  and_inst0__in1;
  wire  and_inst0__out;
  corebit_and and_inst0(
    .in0(and_inst0__in0),
    .in1(and_inst0__in1),
    .out(and_inst0__out)
  );

  // Instancing generated Module: coreir.const(width:8)
  wire [7:0] const_10_8__out;
  coreir_const #(.value(8'h0a),.width(8)) const_10_8(
    .out(const_10_8__out)
  );

  // Instancing generated Module: coreir.eq(width:8)
  wire [7:0] coreir_eq_8_inst0__in0;
  wire [7:0] coreir_eq_8_inst0__in1;
  wire  coreir_eq_8_inst0__out;
  coreir_eq #(.width(8)) coreir_eq_8_inst0(
    .in0(coreir_eq_8_inst0__in0),
    .in1(coreir_eq_8_inst0__in1),
    .out(coreir_eq_8_inst0__out)
  );

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET = reset;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE = and_inst0__out;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK = clk;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I[0] = config_data[0];

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I[1] = config_data[1];

  assign O[1:0] = Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O[1:0];

  assign and_inst0__in0 = coreir_eq_8_inst0__out;

  assign and_inst0__in1 = config_en;

  assign coreir_eq_8_inst0__in1[7:0] = const_10_8__out[7:0];

  assign coreir_eq_8_inst0__in0[7:0] = config_addr[7:0];


endmodule  // ConfigRegister_2_8_32_10

module ConfigRegister_2_8_32_0 (
  output [1:0] O,
  input  clk,
  input [7:0] config_addr,
  input [31:0] config_data,
  input  config_en,
  input  reset
);


  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK;
  wire [1:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I;
  wire [1:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O;
  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2 Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0(
    .ASYNCRESET(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET),
    .CE(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE),
    .CLK(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK),
    .I(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O)
  );

  wire  and_inst0__in0;
  wire  and_inst0__in1;
  wire  and_inst0__out;
  corebit_and and_inst0(
    .in0(and_inst0__in0),
    .in1(and_inst0__in1),
    .out(and_inst0__out)
  );

  // Instancing generated Module: coreir.const(width:8)
  wire [7:0] const_0_8__out;
  coreir_const #(.value(8'h00),.width(8)) const_0_8(
    .out(const_0_8__out)
  );

  // Instancing generated Module: coreir.eq(width:8)
  wire [7:0] coreir_eq_8_inst0__in0;
  wire [7:0] coreir_eq_8_inst0__in1;
  wire  coreir_eq_8_inst0__out;
  coreir_eq #(.width(8)) coreir_eq_8_inst0(
    .in0(coreir_eq_8_inst0__in0),
    .in1(coreir_eq_8_inst0__in1),
    .out(coreir_eq_8_inst0__out)
  );

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__ASYNCRESET = reset;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CE = and_inst0__out;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__CLK = clk;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I[0] = config_data[0];

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__I[1] = config_data[1];

  assign O[1:0] = Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_2_inst0__O[1:0];

  assign and_inst0__in0 = coreir_eq_8_inst0__out;

  assign and_inst0__in1 = config_en;

  assign coreir_eq_8_inst0__in1[7:0] = const_0_8__out[7:0];

  assign coreir_eq_8_inst0__in0[7:0] = config_addr[7:0];


endmodule  // ConfigRegister_2_8_32_0

module ConfigRegister_1_8_32_9 (
  output [0:0] O,
  input  clk,
  input [7:0] config_addr,
  input [31:0] config_data,
  input  config_en,
  input  reset
);


  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__ASYNCRESET;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CE;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CLK;
  wire [0:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__I;
  wire [0:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__O;
  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1 Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0(
    .ASYNCRESET(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__ASYNCRESET),
    .CE(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CE),
    .CLK(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CLK),
    .I(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__I),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__O)
  );

  wire  and_inst0__in0;
  wire  and_inst0__in1;
  wire  and_inst0__out;
  corebit_and and_inst0(
    .in0(and_inst0__in0),
    .in1(and_inst0__in1),
    .out(and_inst0__out)
  );

  // Instancing generated Module: coreir.const(width:8)
  wire [7:0] const_9_8__out;
  coreir_const #(.value(8'h09),.width(8)) const_9_8(
    .out(const_9_8__out)
  );

  // Instancing generated Module: coreir.eq(width:8)
  wire [7:0] coreir_eq_8_inst0__in0;
  wire [7:0] coreir_eq_8_inst0__in1;
  wire  coreir_eq_8_inst0__out;
  coreir_eq #(.width(8)) coreir_eq_8_inst0(
    .in0(coreir_eq_8_inst0__in0),
    .in1(coreir_eq_8_inst0__in1),
    .out(coreir_eq_8_inst0__out)
  );

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__ASYNCRESET = reset;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CE = and_inst0__out;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CLK = clk;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__I[0] = config_data[0];

  assign O[0:0] = Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__O[0:0];

  assign and_inst0__in0 = coreir_eq_8_inst0__out;

  assign and_inst0__in1 = config_en;

  assign coreir_eq_8_inst0__in1[7:0] = const_9_8__out[7:0];

  assign coreir_eq_8_inst0__in0[7:0] = config_addr[7:0];


endmodule  // ConfigRegister_1_8_32_9

module ConfigRegister_1_8_32_79 (
  output [0:0] O,
  input  clk,
  input [7:0] config_addr,
  input [31:0] config_data,
  input  config_en,
  input  reset
);


  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__ASYNCRESET;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CE;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CLK;
  wire [0:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__I;
  wire [0:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__O;
  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1 Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0(
    .ASYNCRESET(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__ASYNCRESET),
    .CE(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CE),
    .CLK(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CLK),
    .I(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__I),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__O)
  );

  wire  and_inst0__in0;
  wire  and_inst0__in1;
  wire  and_inst0__out;
  corebit_and and_inst0(
    .in0(and_inst0__in0),
    .in1(and_inst0__in1),
    .out(and_inst0__out)
  );

  // Instancing generated Module: coreir.const(width:8)
  wire [7:0] const_79_8__out;
  coreir_const #(.value(8'h4f),.width(8)) const_79_8(
    .out(const_79_8__out)
  );

  // Instancing generated Module: coreir.eq(width:8)
  wire [7:0] coreir_eq_8_inst0__in0;
  wire [7:0] coreir_eq_8_inst0__in1;
  wire  coreir_eq_8_inst0__out;
  coreir_eq #(.width(8)) coreir_eq_8_inst0(
    .in0(coreir_eq_8_inst0__in0),
    .in1(coreir_eq_8_inst0__in1),
    .out(coreir_eq_8_inst0__out)
  );

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__ASYNCRESET = reset;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CE = and_inst0__out;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CLK = clk;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__I[0] = config_data[0];

  assign O[0:0] = Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__O[0:0];

  assign and_inst0__in0 = coreir_eq_8_inst0__out;

  assign and_inst0__in1 = config_en;

  assign coreir_eq_8_inst0__in1[7:0] = const_79_8__out[7:0];

  assign coreir_eq_8_inst0__in0[7:0] = config_addr[7:0];


endmodule  // ConfigRegister_1_8_32_79

module ConfigRegister_1_8_32_77 (
  output [0:0] O,
  input  clk,
  input [7:0] config_addr,
  input [31:0] config_data,
  input  config_en,
  input  reset
);


  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__ASYNCRESET;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CE;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CLK;
  wire [0:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__I;
  wire [0:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__O;
  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1 Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0(
    .ASYNCRESET(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__ASYNCRESET),
    .CE(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CE),
    .CLK(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CLK),
    .I(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__I),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__O)
  );

  wire  and_inst0__in0;
  wire  and_inst0__in1;
  wire  and_inst0__out;
  corebit_and and_inst0(
    .in0(and_inst0__in0),
    .in1(and_inst0__in1),
    .out(and_inst0__out)
  );

  // Instancing generated Module: coreir.const(width:8)
  wire [7:0] const_77_8__out;
  coreir_const #(.value(8'h4d),.width(8)) const_77_8(
    .out(const_77_8__out)
  );

  // Instancing generated Module: coreir.eq(width:8)
  wire [7:0] coreir_eq_8_inst0__in0;
  wire [7:0] coreir_eq_8_inst0__in1;
  wire  coreir_eq_8_inst0__out;
  coreir_eq #(.width(8)) coreir_eq_8_inst0(
    .in0(coreir_eq_8_inst0__in0),
    .in1(coreir_eq_8_inst0__in1),
    .out(coreir_eq_8_inst0__out)
  );

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__ASYNCRESET = reset;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CE = and_inst0__out;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CLK = clk;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__I[0] = config_data[0];

  assign O[0:0] = Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__O[0:0];

  assign and_inst0__in0 = coreir_eq_8_inst0__out;

  assign and_inst0__in1 = config_en;

  assign coreir_eq_8_inst0__in1[7:0] = const_77_8__out[7:0];

  assign coreir_eq_8_inst0__in0[7:0] = config_addr[7:0];


endmodule  // ConfigRegister_1_8_32_77

module ConfigRegister_1_8_32_75 (
  output [0:0] O,
  input  clk,
  input [7:0] config_addr,
  input [31:0] config_data,
  input  config_en,
  input  reset
);


  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__ASYNCRESET;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CE;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CLK;
  wire [0:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__I;
  wire [0:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__O;
  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1 Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0(
    .ASYNCRESET(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__ASYNCRESET),
    .CE(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CE),
    .CLK(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CLK),
    .I(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__I),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__O)
  );

  wire  and_inst0__in0;
  wire  and_inst0__in1;
  wire  and_inst0__out;
  corebit_and and_inst0(
    .in0(and_inst0__in0),
    .in1(and_inst0__in1),
    .out(and_inst0__out)
  );

  // Instancing generated Module: coreir.const(width:8)
  wire [7:0] const_75_8__out;
  coreir_const #(.value(8'h4b),.width(8)) const_75_8(
    .out(const_75_8__out)
  );

  // Instancing generated Module: coreir.eq(width:8)
  wire [7:0] coreir_eq_8_inst0__in0;
  wire [7:0] coreir_eq_8_inst0__in1;
  wire  coreir_eq_8_inst0__out;
  coreir_eq #(.width(8)) coreir_eq_8_inst0(
    .in0(coreir_eq_8_inst0__in0),
    .in1(coreir_eq_8_inst0__in1),
    .out(coreir_eq_8_inst0__out)
  );

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__ASYNCRESET = reset;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CE = and_inst0__out;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CLK = clk;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__I[0] = config_data[0];

  assign O[0:0] = Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__O[0:0];

  assign and_inst0__in0 = coreir_eq_8_inst0__out;

  assign and_inst0__in1 = config_en;

  assign coreir_eq_8_inst0__in1[7:0] = const_75_8__out[7:0];

  assign coreir_eq_8_inst0__in0[7:0] = config_addr[7:0];


endmodule  // ConfigRegister_1_8_32_75

module ConfigRegister_1_8_32_73 (
  output [0:0] O,
  input  clk,
  input [7:0] config_addr,
  input [31:0] config_data,
  input  config_en,
  input  reset
);


  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__ASYNCRESET;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CE;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CLK;
  wire [0:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__I;
  wire [0:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__O;
  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1 Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0(
    .ASYNCRESET(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__ASYNCRESET),
    .CE(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CE),
    .CLK(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CLK),
    .I(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__I),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__O)
  );

  wire  and_inst0__in0;
  wire  and_inst0__in1;
  wire  and_inst0__out;
  corebit_and and_inst0(
    .in0(and_inst0__in0),
    .in1(and_inst0__in1),
    .out(and_inst0__out)
  );

  // Instancing generated Module: coreir.const(width:8)
  wire [7:0] const_73_8__out;
  coreir_const #(.value(8'h49),.width(8)) const_73_8(
    .out(const_73_8__out)
  );

  // Instancing generated Module: coreir.eq(width:8)
  wire [7:0] coreir_eq_8_inst0__in0;
  wire [7:0] coreir_eq_8_inst0__in1;
  wire  coreir_eq_8_inst0__out;
  coreir_eq #(.width(8)) coreir_eq_8_inst0(
    .in0(coreir_eq_8_inst0__in0),
    .in1(coreir_eq_8_inst0__in1),
    .out(coreir_eq_8_inst0__out)
  );

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__ASYNCRESET = reset;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CE = and_inst0__out;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CLK = clk;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__I[0] = config_data[0];

  assign O[0:0] = Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__O[0:0];

  assign and_inst0__in0 = coreir_eq_8_inst0__out;

  assign and_inst0__in1 = config_en;

  assign coreir_eq_8_inst0__in1[7:0] = const_73_8__out[7:0];

  assign coreir_eq_8_inst0__in0[7:0] = config_addr[7:0];


endmodule  // ConfigRegister_1_8_32_73

module ConfigRegister_1_8_32_71 (
  output [0:0] O,
  input  clk,
  input [7:0] config_addr,
  input [31:0] config_data,
  input  config_en,
  input  reset
);


  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__ASYNCRESET;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CE;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CLK;
  wire [0:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__I;
  wire [0:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__O;
  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1 Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0(
    .ASYNCRESET(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__ASYNCRESET),
    .CE(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CE),
    .CLK(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CLK),
    .I(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__I),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__O)
  );

  wire  and_inst0__in0;
  wire  and_inst0__in1;
  wire  and_inst0__out;
  corebit_and and_inst0(
    .in0(and_inst0__in0),
    .in1(and_inst0__in1),
    .out(and_inst0__out)
  );

  // Instancing generated Module: coreir.const(width:8)
  wire [7:0] const_71_8__out;
  coreir_const #(.value(8'h47),.width(8)) const_71_8(
    .out(const_71_8__out)
  );

  // Instancing generated Module: coreir.eq(width:8)
  wire [7:0] coreir_eq_8_inst0__in0;
  wire [7:0] coreir_eq_8_inst0__in1;
  wire  coreir_eq_8_inst0__out;
  coreir_eq #(.width(8)) coreir_eq_8_inst0(
    .in0(coreir_eq_8_inst0__in0),
    .in1(coreir_eq_8_inst0__in1),
    .out(coreir_eq_8_inst0__out)
  );

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__ASYNCRESET = reset;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CE = and_inst0__out;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CLK = clk;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__I[0] = config_data[0];

  assign O[0:0] = Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__O[0:0];

  assign and_inst0__in0 = coreir_eq_8_inst0__out;

  assign and_inst0__in1 = config_en;

  assign coreir_eq_8_inst0__in1[7:0] = const_71_8__out[7:0];

  assign coreir_eq_8_inst0__in0[7:0] = config_addr[7:0];


endmodule  // ConfigRegister_1_8_32_71

module ConfigRegister_1_8_32_7 (
  output [0:0] O,
  input  clk,
  input [7:0] config_addr,
  input [31:0] config_data,
  input  config_en,
  input  reset
);


  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__ASYNCRESET;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CE;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CLK;
  wire [0:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__I;
  wire [0:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__O;
  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1 Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0(
    .ASYNCRESET(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__ASYNCRESET),
    .CE(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CE),
    .CLK(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CLK),
    .I(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__I),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__O)
  );

  wire  and_inst0__in0;
  wire  and_inst0__in1;
  wire  and_inst0__out;
  corebit_and and_inst0(
    .in0(and_inst0__in0),
    .in1(and_inst0__in1),
    .out(and_inst0__out)
  );

  // Instancing generated Module: coreir.const(width:8)
  wire [7:0] const_7_8__out;
  coreir_const #(.value(8'h07),.width(8)) const_7_8(
    .out(const_7_8__out)
  );

  // Instancing generated Module: coreir.eq(width:8)
  wire [7:0] coreir_eq_8_inst0__in0;
  wire [7:0] coreir_eq_8_inst0__in1;
  wire  coreir_eq_8_inst0__out;
  coreir_eq #(.width(8)) coreir_eq_8_inst0(
    .in0(coreir_eq_8_inst0__in0),
    .in1(coreir_eq_8_inst0__in1),
    .out(coreir_eq_8_inst0__out)
  );

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__ASYNCRESET = reset;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CE = and_inst0__out;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CLK = clk;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__I[0] = config_data[0];

  assign O[0:0] = Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__O[0:0];

  assign and_inst0__in0 = coreir_eq_8_inst0__out;

  assign and_inst0__in1 = config_en;

  assign coreir_eq_8_inst0__in1[7:0] = const_7_8__out[7:0];

  assign coreir_eq_8_inst0__in0[7:0] = config_addr[7:0];


endmodule  // ConfigRegister_1_8_32_7

module ConfigRegister_1_8_32_69 (
  output [0:0] O,
  input  clk,
  input [7:0] config_addr,
  input [31:0] config_data,
  input  config_en,
  input  reset
);


  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__ASYNCRESET;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CE;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CLK;
  wire [0:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__I;
  wire [0:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__O;
  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1 Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0(
    .ASYNCRESET(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__ASYNCRESET),
    .CE(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CE),
    .CLK(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CLK),
    .I(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__I),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__O)
  );

  wire  and_inst0__in0;
  wire  and_inst0__in1;
  wire  and_inst0__out;
  corebit_and and_inst0(
    .in0(and_inst0__in0),
    .in1(and_inst0__in1),
    .out(and_inst0__out)
  );

  // Instancing generated Module: coreir.const(width:8)
  wire [7:0] const_69_8__out;
  coreir_const #(.value(8'h45),.width(8)) const_69_8(
    .out(const_69_8__out)
  );

  // Instancing generated Module: coreir.eq(width:8)
  wire [7:0] coreir_eq_8_inst0__in0;
  wire [7:0] coreir_eq_8_inst0__in1;
  wire  coreir_eq_8_inst0__out;
  coreir_eq #(.width(8)) coreir_eq_8_inst0(
    .in0(coreir_eq_8_inst0__in0),
    .in1(coreir_eq_8_inst0__in1),
    .out(coreir_eq_8_inst0__out)
  );

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__ASYNCRESET = reset;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CE = and_inst0__out;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CLK = clk;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__I[0] = config_data[0];

  assign O[0:0] = Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__O[0:0];

  assign and_inst0__in0 = coreir_eq_8_inst0__out;

  assign and_inst0__in1 = config_en;

  assign coreir_eq_8_inst0__in1[7:0] = const_69_8__out[7:0];

  assign coreir_eq_8_inst0__in0[7:0] = config_addr[7:0];


endmodule  // ConfigRegister_1_8_32_69

module ConfigRegister_1_8_32_67 (
  output [0:0] O,
  input  clk,
  input [7:0] config_addr,
  input [31:0] config_data,
  input  config_en,
  input  reset
);


  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__ASYNCRESET;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CE;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CLK;
  wire [0:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__I;
  wire [0:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__O;
  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1 Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0(
    .ASYNCRESET(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__ASYNCRESET),
    .CE(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CE),
    .CLK(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CLK),
    .I(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__I),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__O)
  );

  wire  and_inst0__in0;
  wire  and_inst0__in1;
  wire  and_inst0__out;
  corebit_and and_inst0(
    .in0(and_inst0__in0),
    .in1(and_inst0__in1),
    .out(and_inst0__out)
  );

  // Instancing generated Module: coreir.const(width:8)
  wire [7:0] const_67_8__out;
  coreir_const #(.value(8'h43),.width(8)) const_67_8(
    .out(const_67_8__out)
  );

  // Instancing generated Module: coreir.eq(width:8)
  wire [7:0] coreir_eq_8_inst0__in0;
  wire [7:0] coreir_eq_8_inst0__in1;
  wire  coreir_eq_8_inst0__out;
  coreir_eq #(.width(8)) coreir_eq_8_inst0(
    .in0(coreir_eq_8_inst0__in0),
    .in1(coreir_eq_8_inst0__in1),
    .out(coreir_eq_8_inst0__out)
  );

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__ASYNCRESET = reset;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CE = and_inst0__out;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CLK = clk;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__I[0] = config_data[0];

  assign O[0:0] = Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__O[0:0];

  assign and_inst0__in0 = coreir_eq_8_inst0__out;

  assign and_inst0__in1 = config_en;

  assign coreir_eq_8_inst0__in1[7:0] = const_67_8__out[7:0];

  assign coreir_eq_8_inst0__in0[7:0] = config_addr[7:0];


endmodule  // ConfigRegister_1_8_32_67

module ConfigRegister_1_8_32_65 (
  output [0:0] O,
  input  clk,
  input [7:0] config_addr,
  input [31:0] config_data,
  input  config_en,
  input  reset
);


  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__ASYNCRESET;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CE;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CLK;
  wire [0:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__I;
  wire [0:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__O;
  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1 Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0(
    .ASYNCRESET(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__ASYNCRESET),
    .CE(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CE),
    .CLK(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CLK),
    .I(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__I),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__O)
  );

  wire  and_inst0__in0;
  wire  and_inst0__in1;
  wire  and_inst0__out;
  corebit_and and_inst0(
    .in0(and_inst0__in0),
    .in1(and_inst0__in1),
    .out(and_inst0__out)
  );

  // Instancing generated Module: coreir.const(width:8)
  wire [7:0] const_65_8__out;
  coreir_const #(.value(8'h41),.width(8)) const_65_8(
    .out(const_65_8__out)
  );

  // Instancing generated Module: coreir.eq(width:8)
  wire [7:0] coreir_eq_8_inst0__in0;
  wire [7:0] coreir_eq_8_inst0__in1;
  wire  coreir_eq_8_inst0__out;
  coreir_eq #(.width(8)) coreir_eq_8_inst0(
    .in0(coreir_eq_8_inst0__in0),
    .in1(coreir_eq_8_inst0__in1),
    .out(coreir_eq_8_inst0__out)
  );

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__ASYNCRESET = reset;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CE = and_inst0__out;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CLK = clk;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__I[0] = config_data[0];

  assign O[0:0] = Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__O[0:0];

  assign and_inst0__in0 = coreir_eq_8_inst0__out;

  assign and_inst0__in1 = config_en;

  assign coreir_eq_8_inst0__in1[7:0] = const_65_8__out[7:0];

  assign coreir_eq_8_inst0__in0[7:0] = config_addr[7:0];


endmodule  // ConfigRegister_1_8_32_65

module ConfigRegister_1_8_32_63 (
  output [0:0] O,
  input  clk,
  input [7:0] config_addr,
  input [31:0] config_data,
  input  config_en,
  input  reset
);


  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__ASYNCRESET;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CE;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CLK;
  wire [0:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__I;
  wire [0:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__O;
  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1 Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0(
    .ASYNCRESET(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__ASYNCRESET),
    .CE(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CE),
    .CLK(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CLK),
    .I(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__I),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__O)
  );

  wire  and_inst0__in0;
  wire  and_inst0__in1;
  wire  and_inst0__out;
  corebit_and and_inst0(
    .in0(and_inst0__in0),
    .in1(and_inst0__in1),
    .out(and_inst0__out)
  );

  // Instancing generated Module: coreir.const(width:8)
  wire [7:0] const_63_8__out;
  coreir_const #(.value(8'h3f),.width(8)) const_63_8(
    .out(const_63_8__out)
  );

  // Instancing generated Module: coreir.eq(width:8)
  wire [7:0] coreir_eq_8_inst0__in0;
  wire [7:0] coreir_eq_8_inst0__in1;
  wire  coreir_eq_8_inst0__out;
  coreir_eq #(.width(8)) coreir_eq_8_inst0(
    .in0(coreir_eq_8_inst0__in0),
    .in1(coreir_eq_8_inst0__in1),
    .out(coreir_eq_8_inst0__out)
  );

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__ASYNCRESET = reset;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CE = and_inst0__out;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CLK = clk;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__I[0] = config_data[0];

  assign O[0:0] = Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__O[0:0];

  assign and_inst0__in0 = coreir_eq_8_inst0__out;

  assign and_inst0__in1 = config_en;

  assign coreir_eq_8_inst0__in1[7:0] = const_63_8__out[7:0];

  assign coreir_eq_8_inst0__in0[7:0] = config_addr[7:0];


endmodule  // ConfigRegister_1_8_32_63

module ConfigRegister_1_8_32_61 (
  output [0:0] O,
  input  clk,
  input [7:0] config_addr,
  input [31:0] config_data,
  input  config_en,
  input  reset
);


  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__ASYNCRESET;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CE;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CLK;
  wire [0:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__I;
  wire [0:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__O;
  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1 Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0(
    .ASYNCRESET(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__ASYNCRESET),
    .CE(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CE),
    .CLK(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CLK),
    .I(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__I),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__O)
  );

  wire  and_inst0__in0;
  wire  and_inst0__in1;
  wire  and_inst0__out;
  corebit_and and_inst0(
    .in0(and_inst0__in0),
    .in1(and_inst0__in1),
    .out(and_inst0__out)
  );

  // Instancing generated Module: coreir.const(width:8)
  wire [7:0] const_61_8__out;
  coreir_const #(.value(8'h3d),.width(8)) const_61_8(
    .out(const_61_8__out)
  );

  // Instancing generated Module: coreir.eq(width:8)
  wire [7:0] coreir_eq_8_inst0__in0;
  wire [7:0] coreir_eq_8_inst0__in1;
  wire  coreir_eq_8_inst0__out;
  coreir_eq #(.width(8)) coreir_eq_8_inst0(
    .in0(coreir_eq_8_inst0__in0),
    .in1(coreir_eq_8_inst0__in1),
    .out(coreir_eq_8_inst0__out)
  );

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__ASYNCRESET = reset;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CE = and_inst0__out;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CLK = clk;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__I[0] = config_data[0];

  assign O[0:0] = Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__O[0:0];

  assign and_inst0__in0 = coreir_eq_8_inst0__out;

  assign and_inst0__in1 = config_en;

  assign coreir_eq_8_inst0__in1[7:0] = const_61_8__out[7:0];

  assign coreir_eq_8_inst0__in0[7:0] = config_addr[7:0];


endmodule  // ConfigRegister_1_8_32_61

module ConfigRegister_1_8_32_59 (
  output [0:0] O,
  input  clk,
  input [7:0] config_addr,
  input [31:0] config_data,
  input  config_en,
  input  reset
);


  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__ASYNCRESET;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CE;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CLK;
  wire [0:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__I;
  wire [0:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__O;
  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1 Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0(
    .ASYNCRESET(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__ASYNCRESET),
    .CE(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CE),
    .CLK(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CLK),
    .I(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__I),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__O)
  );

  wire  and_inst0__in0;
  wire  and_inst0__in1;
  wire  and_inst0__out;
  corebit_and and_inst0(
    .in0(and_inst0__in0),
    .in1(and_inst0__in1),
    .out(and_inst0__out)
  );

  // Instancing generated Module: coreir.const(width:8)
  wire [7:0] const_59_8__out;
  coreir_const #(.value(8'h3b),.width(8)) const_59_8(
    .out(const_59_8__out)
  );

  // Instancing generated Module: coreir.eq(width:8)
  wire [7:0] coreir_eq_8_inst0__in0;
  wire [7:0] coreir_eq_8_inst0__in1;
  wire  coreir_eq_8_inst0__out;
  coreir_eq #(.width(8)) coreir_eq_8_inst0(
    .in0(coreir_eq_8_inst0__in0),
    .in1(coreir_eq_8_inst0__in1),
    .out(coreir_eq_8_inst0__out)
  );

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__ASYNCRESET = reset;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CE = and_inst0__out;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CLK = clk;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__I[0] = config_data[0];

  assign O[0:0] = Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__O[0:0];

  assign and_inst0__in0 = coreir_eq_8_inst0__out;

  assign and_inst0__in1 = config_en;

  assign coreir_eq_8_inst0__in1[7:0] = const_59_8__out[7:0];

  assign coreir_eq_8_inst0__in0[7:0] = config_addr[7:0];


endmodule  // ConfigRegister_1_8_32_59

module ConfigRegister_1_8_32_57 (
  output [0:0] O,
  input  clk,
  input [7:0] config_addr,
  input [31:0] config_data,
  input  config_en,
  input  reset
);


  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__ASYNCRESET;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CE;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CLK;
  wire [0:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__I;
  wire [0:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__O;
  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1 Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0(
    .ASYNCRESET(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__ASYNCRESET),
    .CE(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CE),
    .CLK(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CLK),
    .I(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__I),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__O)
  );

  wire  and_inst0__in0;
  wire  and_inst0__in1;
  wire  and_inst0__out;
  corebit_and and_inst0(
    .in0(and_inst0__in0),
    .in1(and_inst0__in1),
    .out(and_inst0__out)
  );

  // Instancing generated Module: coreir.const(width:8)
  wire [7:0] const_57_8__out;
  coreir_const #(.value(8'h39),.width(8)) const_57_8(
    .out(const_57_8__out)
  );

  // Instancing generated Module: coreir.eq(width:8)
  wire [7:0] coreir_eq_8_inst0__in0;
  wire [7:0] coreir_eq_8_inst0__in1;
  wire  coreir_eq_8_inst0__out;
  coreir_eq #(.width(8)) coreir_eq_8_inst0(
    .in0(coreir_eq_8_inst0__in0),
    .in1(coreir_eq_8_inst0__in1),
    .out(coreir_eq_8_inst0__out)
  );

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__ASYNCRESET = reset;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CE = and_inst0__out;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CLK = clk;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__I[0] = config_data[0];

  assign O[0:0] = Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__O[0:0];

  assign and_inst0__in0 = coreir_eq_8_inst0__out;

  assign and_inst0__in1 = config_en;

  assign coreir_eq_8_inst0__in1[7:0] = const_57_8__out[7:0];

  assign coreir_eq_8_inst0__in0[7:0] = config_addr[7:0];


endmodule  // ConfigRegister_1_8_32_57

module ConfigRegister_1_8_32_55 (
  output [0:0] O,
  input  clk,
  input [7:0] config_addr,
  input [31:0] config_data,
  input  config_en,
  input  reset
);


  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__ASYNCRESET;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CE;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CLK;
  wire [0:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__I;
  wire [0:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__O;
  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1 Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0(
    .ASYNCRESET(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__ASYNCRESET),
    .CE(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CE),
    .CLK(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CLK),
    .I(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__I),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__O)
  );

  wire  and_inst0__in0;
  wire  and_inst0__in1;
  wire  and_inst0__out;
  corebit_and and_inst0(
    .in0(and_inst0__in0),
    .in1(and_inst0__in1),
    .out(and_inst0__out)
  );

  // Instancing generated Module: coreir.const(width:8)
  wire [7:0] const_55_8__out;
  coreir_const #(.value(8'h37),.width(8)) const_55_8(
    .out(const_55_8__out)
  );

  // Instancing generated Module: coreir.eq(width:8)
  wire [7:0] coreir_eq_8_inst0__in0;
  wire [7:0] coreir_eq_8_inst0__in1;
  wire  coreir_eq_8_inst0__out;
  coreir_eq #(.width(8)) coreir_eq_8_inst0(
    .in0(coreir_eq_8_inst0__in0),
    .in1(coreir_eq_8_inst0__in1),
    .out(coreir_eq_8_inst0__out)
  );

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__ASYNCRESET = reset;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CE = and_inst0__out;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CLK = clk;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__I[0] = config_data[0];

  assign O[0:0] = Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__O[0:0];

  assign and_inst0__in0 = coreir_eq_8_inst0__out;

  assign and_inst0__in1 = config_en;

  assign coreir_eq_8_inst0__in1[7:0] = const_55_8__out[7:0];

  assign coreir_eq_8_inst0__in0[7:0] = config_addr[7:0];


endmodule  // ConfigRegister_1_8_32_55

module ConfigRegister_1_8_32_53 (
  output [0:0] O,
  input  clk,
  input [7:0] config_addr,
  input [31:0] config_data,
  input  config_en,
  input  reset
);


  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__ASYNCRESET;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CE;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CLK;
  wire [0:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__I;
  wire [0:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__O;
  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1 Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0(
    .ASYNCRESET(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__ASYNCRESET),
    .CE(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CE),
    .CLK(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CLK),
    .I(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__I),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__O)
  );

  wire  and_inst0__in0;
  wire  and_inst0__in1;
  wire  and_inst0__out;
  corebit_and and_inst0(
    .in0(and_inst0__in0),
    .in1(and_inst0__in1),
    .out(and_inst0__out)
  );

  // Instancing generated Module: coreir.const(width:8)
  wire [7:0] const_53_8__out;
  coreir_const #(.value(8'h35),.width(8)) const_53_8(
    .out(const_53_8__out)
  );

  // Instancing generated Module: coreir.eq(width:8)
  wire [7:0] coreir_eq_8_inst0__in0;
  wire [7:0] coreir_eq_8_inst0__in1;
  wire  coreir_eq_8_inst0__out;
  coreir_eq #(.width(8)) coreir_eq_8_inst0(
    .in0(coreir_eq_8_inst0__in0),
    .in1(coreir_eq_8_inst0__in1),
    .out(coreir_eq_8_inst0__out)
  );

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__ASYNCRESET = reset;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CE = and_inst0__out;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CLK = clk;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__I[0] = config_data[0];

  assign O[0:0] = Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__O[0:0];

  assign and_inst0__in0 = coreir_eq_8_inst0__out;

  assign and_inst0__in1 = config_en;

  assign coreir_eq_8_inst0__in1[7:0] = const_53_8__out[7:0];

  assign coreir_eq_8_inst0__in0[7:0] = config_addr[7:0];


endmodule  // ConfigRegister_1_8_32_53

module ConfigRegister_1_8_32_51 (
  output [0:0] O,
  input  clk,
  input [7:0] config_addr,
  input [31:0] config_data,
  input  config_en,
  input  reset
);


  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__ASYNCRESET;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CE;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CLK;
  wire [0:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__I;
  wire [0:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__O;
  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1 Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0(
    .ASYNCRESET(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__ASYNCRESET),
    .CE(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CE),
    .CLK(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CLK),
    .I(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__I),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__O)
  );

  wire  and_inst0__in0;
  wire  and_inst0__in1;
  wire  and_inst0__out;
  corebit_and and_inst0(
    .in0(and_inst0__in0),
    .in1(and_inst0__in1),
    .out(and_inst0__out)
  );

  // Instancing generated Module: coreir.const(width:8)
  wire [7:0] const_51_8__out;
  coreir_const #(.value(8'h33),.width(8)) const_51_8(
    .out(const_51_8__out)
  );

  // Instancing generated Module: coreir.eq(width:8)
  wire [7:0] coreir_eq_8_inst0__in0;
  wire [7:0] coreir_eq_8_inst0__in1;
  wire  coreir_eq_8_inst0__out;
  coreir_eq #(.width(8)) coreir_eq_8_inst0(
    .in0(coreir_eq_8_inst0__in0),
    .in1(coreir_eq_8_inst0__in1),
    .out(coreir_eq_8_inst0__out)
  );

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__ASYNCRESET = reset;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CE = and_inst0__out;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CLK = clk;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__I[0] = config_data[0];

  assign O[0:0] = Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__O[0:0];

  assign and_inst0__in0 = coreir_eq_8_inst0__out;

  assign and_inst0__in1 = config_en;

  assign coreir_eq_8_inst0__in1[7:0] = const_51_8__out[7:0];

  assign coreir_eq_8_inst0__in0[7:0] = config_addr[7:0];


endmodule  // ConfigRegister_1_8_32_51

module ConfigRegister_1_8_32_5 (
  output [0:0] O,
  input  clk,
  input [7:0] config_addr,
  input [31:0] config_data,
  input  config_en,
  input  reset
);


  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__ASYNCRESET;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CE;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CLK;
  wire [0:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__I;
  wire [0:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__O;
  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1 Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0(
    .ASYNCRESET(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__ASYNCRESET),
    .CE(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CE),
    .CLK(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CLK),
    .I(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__I),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__O)
  );

  wire  and_inst0__in0;
  wire  and_inst0__in1;
  wire  and_inst0__out;
  corebit_and and_inst0(
    .in0(and_inst0__in0),
    .in1(and_inst0__in1),
    .out(and_inst0__out)
  );

  // Instancing generated Module: coreir.const(width:8)
  wire [7:0] const_5_8__out;
  coreir_const #(.value(8'h05),.width(8)) const_5_8(
    .out(const_5_8__out)
  );

  // Instancing generated Module: coreir.eq(width:8)
  wire [7:0] coreir_eq_8_inst0__in0;
  wire [7:0] coreir_eq_8_inst0__in1;
  wire  coreir_eq_8_inst0__out;
  coreir_eq #(.width(8)) coreir_eq_8_inst0(
    .in0(coreir_eq_8_inst0__in0),
    .in1(coreir_eq_8_inst0__in1),
    .out(coreir_eq_8_inst0__out)
  );

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__ASYNCRESET = reset;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CE = and_inst0__out;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CLK = clk;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__I[0] = config_data[0];

  assign O[0:0] = Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__O[0:0];

  assign and_inst0__in0 = coreir_eq_8_inst0__out;

  assign and_inst0__in1 = config_en;

  assign coreir_eq_8_inst0__in1[7:0] = const_5_8__out[7:0];

  assign coreir_eq_8_inst0__in0[7:0] = config_addr[7:0];


endmodule  // ConfigRegister_1_8_32_5

module ConfigRegister_1_8_32_49 (
  output [0:0] O,
  input  clk,
  input [7:0] config_addr,
  input [31:0] config_data,
  input  config_en,
  input  reset
);


  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__ASYNCRESET;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CE;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CLK;
  wire [0:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__I;
  wire [0:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__O;
  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1 Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0(
    .ASYNCRESET(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__ASYNCRESET),
    .CE(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CE),
    .CLK(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CLK),
    .I(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__I),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__O)
  );

  wire  and_inst0__in0;
  wire  and_inst0__in1;
  wire  and_inst0__out;
  corebit_and and_inst0(
    .in0(and_inst0__in0),
    .in1(and_inst0__in1),
    .out(and_inst0__out)
  );

  // Instancing generated Module: coreir.const(width:8)
  wire [7:0] const_49_8__out;
  coreir_const #(.value(8'h31),.width(8)) const_49_8(
    .out(const_49_8__out)
  );

  // Instancing generated Module: coreir.eq(width:8)
  wire [7:0] coreir_eq_8_inst0__in0;
  wire [7:0] coreir_eq_8_inst0__in1;
  wire  coreir_eq_8_inst0__out;
  coreir_eq #(.width(8)) coreir_eq_8_inst0(
    .in0(coreir_eq_8_inst0__in0),
    .in1(coreir_eq_8_inst0__in1),
    .out(coreir_eq_8_inst0__out)
  );

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__ASYNCRESET = reset;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CE = and_inst0__out;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CLK = clk;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__I[0] = config_data[0];

  assign O[0:0] = Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__O[0:0];

  assign and_inst0__in0 = coreir_eq_8_inst0__out;

  assign and_inst0__in1 = config_en;

  assign coreir_eq_8_inst0__in1[7:0] = const_49_8__out[7:0];

  assign coreir_eq_8_inst0__in0[7:0] = config_addr[7:0];


endmodule  // ConfigRegister_1_8_32_49

module ConfigRegister_1_8_32_47 (
  output [0:0] O,
  input  clk,
  input [7:0] config_addr,
  input [31:0] config_data,
  input  config_en,
  input  reset
);


  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__ASYNCRESET;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CE;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CLK;
  wire [0:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__I;
  wire [0:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__O;
  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1 Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0(
    .ASYNCRESET(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__ASYNCRESET),
    .CE(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CE),
    .CLK(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CLK),
    .I(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__I),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__O)
  );

  wire  and_inst0__in0;
  wire  and_inst0__in1;
  wire  and_inst0__out;
  corebit_and and_inst0(
    .in0(and_inst0__in0),
    .in1(and_inst0__in1),
    .out(and_inst0__out)
  );

  // Instancing generated Module: coreir.const(width:8)
  wire [7:0] const_47_8__out;
  coreir_const #(.value(8'h2f),.width(8)) const_47_8(
    .out(const_47_8__out)
  );

  // Instancing generated Module: coreir.eq(width:8)
  wire [7:0] coreir_eq_8_inst0__in0;
  wire [7:0] coreir_eq_8_inst0__in1;
  wire  coreir_eq_8_inst0__out;
  coreir_eq #(.width(8)) coreir_eq_8_inst0(
    .in0(coreir_eq_8_inst0__in0),
    .in1(coreir_eq_8_inst0__in1),
    .out(coreir_eq_8_inst0__out)
  );

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__ASYNCRESET = reset;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CE = and_inst0__out;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CLK = clk;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__I[0] = config_data[0];

  assign O[0:0] = Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__O[0:0];

  assign and_inst0__in0 = coreir_eq_8_inst0__out;

  assign and_inst0__in1 = config_en;

  assign coreir_eq_8_inst0__in1[7:0] = const_47_8__out[7:0];

  assign coreir_eq_8_inst0__in0[7:0] = config_addr[7:0];


endmodule  // ConfigRegister_1_8_32_47

module ConfigRegister_1_8_32_45 (
  output [0:0] O,
  input  clk,
  input [7:0] config_addr,
  input [31:0] config_data,
  input  config_en,
  input  reset
);


  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__ASYNCRESET;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CE;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CLK;
  wire [0:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__I;
  wire [0:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__O;
  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1 Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0(
    .ASYNCRESET(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__ASYNCRESET),
    .CE(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CE),
    .CLK(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CLK),
    .I(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__I),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__O)
  );

  wire  and_inst0__in0;
  wire  and_inst0__in1;
  wire  and_inst0__out;
  corebit_and and_inst0(
    .in0(and_inst0__in0),
    .in1(and_inst0__in1),
    .out(and_inst0__out)
  );

  // Instancing generated Module: coreir.const(width:8)
  wire [7:0] const_45_8__out;
  coreir_const #(.value(8'h2d),.width(8)) const_45_8(
    .out(const_45_8__out)
  );

  // Instancing generated Module: coreir.eq(width:8)
  wire [7:0] coreir_eq_8_inst0__in0;
  wire [7:0] coreir_eq_8_inst0__in1;
  wire  coreir_eq_8_inst0__out;
  coreir_eq #(.width(8)) coreir_eq_8_inst0(
    .in0(coreir_eq_8_inst0__in0),
    .in1(coreir_eq_8_inst0__in1),
    .out(coreir_eq_8_inst0__out)
  );

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__ASYNCRESET = reset;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CE = and_inst0__out;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CLK = clk;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__I[0] = config_data[0];

  assign O[0:0] = Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__O[0:0];

  assign and_inst0__in0 = coreir_eq_8_inst0__out;

  assign and_inst0__in1 = config_en;

  assign coreir_eq_8_inst0__in1[7:0] = const_45_8__out[7:0];

  assign coreir_eq_8_inst0__in0[7:0] = config_addr[7:0];


endmodule  // ConfigRegister_1_8_32_45

module ConfigRegister_1_8_32_43 (
  output [0:0] O,
  input  clk,
  input [7:0] config_addr,
  input [31:0] config_data,
  input  config_en,
  input  reset
);


  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__ASYNCRESET;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CE;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CLK;
  wire [0:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__I;
  wire [0:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__O;
  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1 Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0(
    .ASYNCRESET(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__ASYNCRESET),
    .CE(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CE),
    .CLK(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CLK),
    .I(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__I),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__O)
  );

  wire  and_inst0__in0;
  wire  and_inst0__in1;
  wire  and_inst0__out;
  corebit_and and_inst0(
    .in0(and_inst0__in0),
    .in1(and_inst0__in1),
    .out(and_inst0__out)
  );

  // Instancing generated Module: coreir.const(width:8)
  wire [7:0] const_43_8__out;
  coreir_const #(.value(8'h2b),.width(8)) const_43_8(
    .out(const_43_8__out)
  );

  // Instancing generated Module: coreir.eq(width:8)
  wire [7:0] coreir_eq_8_inst0__in0;
  wire [7:0] coreir_eq_8_inst0__in1;
  wire  coreir_eq_8_inst0__out;
  coreir_eq #(.width(8)) coreir_eq_8_inst0(
    .in0(coreir_eq_8_inst0__in0),
    .in1(coreir_eq_8_inst0__in1),
    .out(coreir_eq_8_inst0__out)
  );

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__ASYNCRESET = reset;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CE = and_inst0__out;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CLK = clk;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__I[0] = config_data[0];

  assign O[0:0] = Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__O[0:0];

  assign and_inst0__in0 = coreir_eq_8_inst0__out;

  assign and_inst0__in1 = config_en;

  assign coreir_eq_8_inst0__in1[7:0] = const_43_8__out[7:0];

  assign coreir_eq_8_inst0__in0[7:0] = config_addr[7:0];


endmodule  // ConfigRegister_1_8_32_43

module ConfigRegister_1_8_32_41 (
  output [0:0] O,
  input  clk,
  input [7:0] config_addr,
  input [31:0] config_data,
  input  config_en,
  input  reset
);


  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__ASYNCRESET;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CE;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CLK;
  wire [0:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__I;
  wire [0:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__O;
  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1 Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0(
    .ASYNCRESET(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__ASYNCRESET),
    .CE(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CE),
    .CLK(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CLK),
    .I(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__I),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__O)
  );

  wire  and_inst0__in0;
  wire  and_inst0__in1;
  wire  and_inst0__out;
  corebit_and and_inst0(
    .in0(and_inst0__in0),
    .in1(and_inst0__in1),
    .out(and_inst0__out)
  );

  // Instancing generated Module: coreir.const(width:8)
  wire [7:0] const_41_8__out;
  coreir_const #(.value(8'h29),.width(8)) const_41_8(
    .out(const_41_8__out)
  );

  // Instancing generated Module: coreir.eq(width:8)
  wire [7:0] coreir_eq_8_inst0__in0;
  wire [7:0] coreir_eq_8_inst0__in1;
  wire  coreir_eq_8_inst0__out;
  coreir_eq #(.width(8)) coreir_eq_8_inst0(
    .in0(coreir_eq_8_inst0__in0),
    .in1(coreir_eq_8_inst0__in1),
    .out(coreir_eq_8_inst0__out)
  );

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__ASYNCRESET = reset;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CE = and_inst0__out;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CLK = clk;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__I[0] = config_data[0];

  assign O[0:0] = Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__O[0:0];

  assign and_inst0__in0 = coreir_eq_8_inst0__out;

  assign and_inst0__in1 = config_en;

  assign coreir_eq_8_inst0__in1[7:0] = const_41_8__out[7:0];

  assign coreir_eq_8_inst0__in0[7:0] = config_addr[7:0];


endmodule  // ConfigRegister_1_8_32_41

module ConfigRegister_1_8_32_39 (
  output [0:0] O,
  input  clk,
  input [7:0] config_addr,
  input [31:0] config_data,
  input  config_en,
  input  reset
);


  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__ASYNCRESET;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CE;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CLK;
  wire [0:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__I;
  wire [0:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__O;
  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1 Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0(
    .ASYNCRESET(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__ASYNCRESET),
    .CE(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CE),
    .CLK(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CLK),
    .I(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__I),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__O)
  );

  wire  and_inst0__in0;
  wire  and_inst0__in1;
  wire  and_inst0__out;
  corebit_and and_inst0(
    .in0(and_inst0__in0),
    .in1(and_inst0__in1),
    .out(and_inst0__out)
  );

  // Instancing generated Module: coreir.const(width:8)
  wire [7:0] const_39_8__out;
  coreir_const #(.value(8'h27),.width(8)) const_39_8(
    .out(const_39_8__out)
  );

  // Instancing generated Module: coreir.eq(width:8)
  wire [7:0] coreir_eq_8_inst0__in0;
  wire [7:0] coreir_eq_8_inst0__in1;
  wire  coreir_eq_8_inst0__out;
  coreir_eq #(.width(8)) coreir_eq_8_inst0(
    .in0(coreir_eq_8_inst0__in0),
    .in1(coreir_eq_8_inst0__in1),
    .out(coreir_eq_8_inst0__out)
  );

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__ASYNCRESET = reset;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CE = and_inst0__out;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CLK = clk;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__I[0] = config_data[0];

  assign O[0:0] = Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__O[0:0];

  assign and_inst0__in0 = coreir_eq_8_inst0__out;

  assign and_inst0__in1 = config_en;

  assign coreir_eq_8_inst0__in1[7:0] = const_39_8__out[7:0];

  assign coreir_eq_8_inst0__in0[7:0] = config_addr[7:0];


endmodule  // ConfigRegister_1_8_32_39

module ConfigRegister_1_8_32_37 (
  output [0:0] O,
  input  clk,
  input [7:0] config_addr,
  input [31:0] config_data,
  input  config_en,
  input  reset
);


  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__ASYNCRESET;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CE;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CLK;
  wire [0:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__I;
  wire [0:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__O;
  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1 Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0(
    .ASYNCRESET(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__ASYNCRESET),
    .CE(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CE),
    .CLK(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CLK),
    .I(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__I),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__O)
  );

  wire  and_inst0__in0;
  wire  and_inst0__in1;
  wire  and_inst0__out;
  corebit_and and_inst0(
    .in0(and_inst0__in0),
    .in1(and_inst0__in1),
    .out(and_inst0__out)
  );

  // Instancing generated Module: coreir.const(width:8)
  wire [7:0] const_37_8__out;
  coreir_const #(.value(8'h25),.width(8)) const_37_8(
    .out(const_37_8__out)
  );

  // Instancing generated Module: coreir.eq(width:8)
  wire [7:0] coreir_eq_8_inst0__in0;
  wire [7:0] coreir_eq_8_inst0__in1;
  wire  coreir_eq_8_inst0__out;
  coreir_eq #(.width(8)) coreir_eq_8_inst0(
    .in0(coreir_eq_8_inst0__in0),
    .in1(coreir_eq_8_inst0__in1),
    .out(coreir_eq_8_inst0__out)
  );

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__ASYNCRESET = reset;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CE = and_inst0__out;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CLK = clk;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__I[0] = config_data[0];

  assign O[0:0] = Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__O[0:0];

  assign and_inst0__in0 = coreir_eq_8_inst0__out;

  assign and_inst0__in1 = config_en;

  assign coreir_eq_8_inst0__in1[7:0] = const_37_8__out[7:0];

  assign coreir_eq_8_inst0__in0[7:0] = config_addr[7:0];


endmodule  // ConfigRegister_1_8_32_37

module ConfigRegister_1_8_32_35 (
  output [0:0] O,
  input  clk,
  input [7:0] config_addr,
  input [31:0] config_data,
  input  config_en,
  input  reset
);


  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__ASYNCRESET;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CE;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CLK;
  wire [0:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__I;
  wire [0:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__O;
  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1 Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0(
    .ASYNCRESET(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__ASYNCRESET),
    .CE(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CE),
    .CLK(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CLK),
    .I(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__I),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__O)
  );

  wire  and_inst0__in0;
  wire  and_inst0__in1;
  wire  and_inst0__out;
  corebit_and and_inst0(
    .in0(and_inst0__in0),
    .in1(and_inst0__in1),
    .out(and_inst0__out)
  );

  // Instancing generated Module: coreir.const(width:8)
  wire [7:0] const_35_8__out;
  coreir_const #(.value(8'h23),.width(8)) const_35_8(
    .out(const_35_8__out)
  );

  // Instancing generated Module: coreir.eq(width:8)
  wire [7:0] coreir_eq_8_inst0__in0;
  wire [7:0] coreir_eq_8_inst0__in1;
  wire  coreir_eq_8_inst0__out;
  coreir_eq #(.width(8)) coreir_eq_8_inst0(
    .in0(coreir_eq_8_inst0__in0),
    .in1(coreir_eq_8_inst0__in1),
    .out(coreir_eq_8_inst0__out)
  );

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__ASYNCRESET = reset;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CE = and_inst0__out;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CLK = clk;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__I[0] = config_data[0];

  assign O[0:0] = Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__O[0:0];

  assign and_inst0__in0 = coreir_eq_8_inst0__out;

  assign and_inst0__in1 = config_en;

  assign coreir_eq_8_inst0__in1[7:0] = const_35_8__out[7:0];

  assign coreir_eq_8_inst0__in0[7:0] = config_addr[7:0];


endmodule  // ConfigRegister_1_8_32_35

module ConfigRegister_1_8_32_33 (
  output [0:0] O,
  input  clk,
  input [7:0] config_addr,
  input [31:0] config_data,
  input  config_en,
  input  reset
);


  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__ASYNCRESET;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CE;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CLK;
  wire [0:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__I;
  wire [0:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__O;
  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1 Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0(
    .ASYNCRESET(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__ASYNCRESET),
    .CE(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CE),
    .CLK(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CLK),
    .I(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__I),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__O)
  );

  wire  and_inst0__in0;
  wire  and_inst0__in1;
  wire  and_inst0__out;
  corebit_and and_inst0(
    .in0(and_inst0__in0),
    .in1(and_inst0__in1),
    .out(and_inst0__out)
  );

  // Instancing generated Module: coreir.const(width:8)
  wire [7:0] const_33_8__out;
  coreir_const #(.value(8'h21),.width(8)) const_33_8(
    .out(const_33_8__out)
  );

  // Instancing generated Module: coreir.eq(width:8)
  wire [7:0] coreir_eq_8_inst0__in0;
  wire [7:0] coreir_eq_8_inst0__in1;
  wire  coreir_eq_8_inst0__out;
  coreir_eq #(.width(8)) coreir_eq_8_inst0(
    .in0(coreir_eq_8_inst0__in0),
    .in1(coreir_eq_8_inst0__in1),
    .out(coreir_eq_8_inst0__out)
  );

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__ASYNCRESET = reset;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CE = and_inst0__out;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CLK = clk;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__I[0] = config_data[0];

  assign O[0:0] = Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__O[0:0];

  assign and_inst0__in0 = coreir_eq_8_inst0__out;

  assign and_inst0__in1 = config_en;

  assign coreir_eq_8_inst0__in1[7:0] = const_33_8__out[7:0];

  assign coreir_eq_8_inst0__in0[7:0] = config_addr[7:0];


endmodule  // ConfigRegister_1_8_32_33

module ConfigRegister_1_8_32_31 (
  output [0:0] O,
  input  clk,
  input [7:0] config_addr,
  input [31:0] config_data,
  input  config_en,
  input  reset
);


  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__ASYNCRESET;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CE;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CLK;
  wire [0:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__I;
  wire [0:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__O;
  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1 Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0(
    .ASYNCRESET(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__ASYNCRESET),
    .CE(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CE),
    .CLK(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CLK),
    .I(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__I),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__O)
  );

  wire  and_inst0__in0;
  wire  and_inst0__in1;
  wire  and_inst0__out;
  corebit_and and_inst0(
    .in0(and_inst0__in0),
    .in1(and_inst0__in1),
    .out(and_inst0__out)
  );

  // Instancing generated Module: coreir.const(width:8)
  wire [7:0] const_31_8__out;
  coreir_const #(.value(8'h1f),.width(8)) const_31_8(
    .out(const_31_8__out)
  );

  // Instancing generated Module: coreir.eq(width:8)
  wire [7:0] coreir_eq_8_inst0__in0;
  wire [7:0] coreir_eq_8_inst0__in1;
  wire  coreir_eq_8_inst0__out;
  coreir_eq #(.width(8)) coreir_eq_8_inst0(
    .in0(coreir_eq_8_inst0__in0),
    .in1(coreir_eq_8_inst0__in1),
    .out(coreir_eq_8_inst0__out)
  );

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__ASYNCRESET = reset;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CE = and_inst0__out;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CLK = clk;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__I[0] = config_data[0];

  assign O[0:0] = Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__O[0:0];

  assign and_inst0__in0 = coreir_eq_8_inst0__out;

  assign and_inst0__in1 = config_en;

  assign coreir_eq_8_inst0__in1[7:0] = const_31_8__out[7:0];

  assign coreir_eq_8_inst0__in0[7:0] = config_addr[7:0];


endmodule  // ConfigRegister_1_8_32_31

module ConfigRegister_1_8_32_3 (
  output [0:0] O,
  input  clk,
  input [7:0] config_addr,
  input [31:0] config_data,
  input  config_en,
  input  reset
);


  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__ASYNCRESET;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CE;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CLK;
  wire [0:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__I;
  wire [0:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__O;
  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1 Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0(
    .ASYNCRESET(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__ASYNCRESET),
    .CE(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CE),
    .CLK(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CLK),
    .I(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__I),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__O)
  );

  wire  and_inst0__in0;
  wire  and_inst0__in1;
  wire  and_inst0__out;
  corebit_and and_inst0(
    .in0(and_inst0__in0),
    .in1(and_inst0__in1),
    .out(and_inst0__out)
  );

  // Instancing generated Module: coreir.const(width:8)
  wire [7:0] const_3_8__out;
  coreir_const #(.value(8'h03),.width(8)) const_3_8(
    .out(const_3_8__out)
  );

  // Instancing generated Module: coreir.eq(width:8)
  wire [7:0] coreir_eq_8_inst0__in0;
  wire [7:0] coreir_eq_8_inst0__in1;
  wire  coreir_eq_8_inst0__out;
  coreir_eq #(.width(8)) coreir_eq_8_inst0(
    .in0(coreir_eq_8_inst0__in0),
    .in1(coreir_eq_8_inst0__in1),
    .out(coreir_eq_8_inst0__out)
  );

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__ASYNCRESET = reset;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CE = and_inst0__out;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CLK = clk;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__I[0] = config_data[0];

  assign O[0:0] = Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__O[0:0];

  assign and_inst0__in0 = coreir_eq_8_inst0__out;

  assign and_inst0__in1 = config_en;

  assign coreir_eq_8_inst0__in1[7:0] = const_3_8__out[7:0];

  assign coreir_eq_8_inst0__in0[7:0] = config_addr[7:0];


endmodule  // ConfigRegister_1_8_32_3

module ConfigRegister_1_8_32_29 (
  output [0:0] O,
  input  clk,
  input [7:0] config_addr,
  input [31:0] config_data,
  input  config_en,
  input  reset
);


  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__ASYNCRESET;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CE;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CLK;
  wire [0:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__I;
  wire [0:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__O;
  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1 Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0(
    .ASYNCRESET(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__ASYNCRESET),
    .CE(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CE),
    .CLK(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CLK),
    .I(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__I),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__O)
  );

  wire  and_inst0__in0;
  wire  and_inst0__in1;
  wire  and_inst0__out;
  corebit_and and_inst0(
    .in0(and_inst0__in0),
    .in1(and_inst0__in1),
    .out(and_inst0__out)
  );

  // Instancing generated Module: coreir.const(width:8)
  wire [7:0] const_29_8__out;
  coreir_const #(.value(8'h1d),.width(8)) const_29_8(
    .out(const_29_8__out)
  );

  // Instancing generated Module: coreir.eq(width:8)
  wire [7:0] coreir_eq_8_inst0__in0;
  wire [7:0] coreir_eq_8_inst0__in1;
  wire  coreir_eq_8_inst0__out;
  coreir_eq #(.width(8)) coreir_eq_8_inst0(
    .in0(coreir_eq_8_inst0__in0),
    .in1(coreir_eq_8_inst0__in1),
    .out(coreir_eq_8_inst0__out)
  );

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__ASYNCRESET = reset;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CE = and_inst0__out;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CLK = clk;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__I[0] = config_data[0];

  assign O[0:0] = Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__O[0:0];

  assign and_inst0__in0 = coreir_eq_8_inst0__out;

  assign and_inst0__in1 = config_en;

  assign coreir_eq_8_inst0__in1[7:0] = const_29_8__out[7:0];

  assign coreir_eq_8_inst0__in0[7:0] = config_addr[7:0];


endmodule  // ConfigRegister_1_8_32_29

module ConfigRegister_1_8_32_27 (
  output [0:0] O,
  input  clk,
  input [7:0] config_addr,
  input [31:0] config_data,
  input  config_en,
  input  reset
);


  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__ASYNCRESET;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CE;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CLK;
  wire [0:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__I;
  wire [0:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__O;
  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1 Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0(
    .ASYNCRESET(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__ASYNCRESET),
    .CE(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CE),
    .CLK(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CLK),
    .I(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__I),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__O)
  );

  wire  and_inst0__in0;
  wire  and_inst0__in1;
  wire  and_inst0__out;
  corebit_and and_inst0(
    .in0(and_inst0__in0),
    .in1(and_inst0__in1),
    .out(and_inst0__out)
  );

  // Instancing generated Module: coreir.const(width:8)
  wire [7:0] const_27_8__out;
  coreir_const #(.value(8'h1b),.width(8)) const_27_8(
    .out(const_27_8__out)
  );

  // Instancing generated Module: coreir.eq(width:8)
  wire [7:0] coreir_eq_8_inst0__in0;
  wire [7:0] coreir_eq_8_inst0__in1;
  wire  coreir_eq_8_inst0__out;
  coreir_eq #(.width(8)) coreir_eq_8_inst0(
    .in0(coreir_eq_8_inst0__in0),
    .in1(coreir_eq_8_inst0__in1),
    .out(coreir_eq_8_inst0__out)
  );

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__ASYNCRESET = reset;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CE = and_inst0__out;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CLK = clk;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__I[0] = config_data[0];

  assign O[0:0] = Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__O[0:0];

  assign and_inst0__in0 = coreir_eq_8_inst0__out;

  assign and_inst0__in1 = config_en;

  assign coreir_eq_8_inst0__in1[7:0] = const_27_8__out[7:0];

  assign coreir_eq_8_inst0__in0[7:0] = config_addr[7:0];


endmodule  // ConfigRegister_1_8_32_27

module ConfigRegister_1_8_32_25 (
  output [0:0] O,
  input  clk,
  input [7:0] config_addr,
  input [31:0] config_data,
  input  config_en,
  input  reset
);


  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__ASYNCRESET;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CE;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CLK;
  wire [0:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__I;
  wire [0:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__O;
  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1 Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0(
    .ASYNCRESET(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__ASYNCRESET),
    .CE(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CE),
    .CLK(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CLK),
    .I(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__I),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__O)
  );

  wire  and_inst0__in0;
  wire  and_inst0__in1;
  wire  and_inst0__out;
  corebit_and and_inst0(
    .in0(and_inst0__in0),
    .in1(and_inst0__in1),
    .out(and_inst0__out)
  );

  // Instancing generated Module: coreir.const(width:8)
  wire [7:0] const_25_8__out;
  coreir_const #(.value(8'h19),.width(8)) const_25_8(
    .out(const_25_8__out)
  );

  // Instancing generated Module: coreir.eq(width:8)
  wire [7:0] coreir_eq_8_inst0__in0;
  wire [7:0] coreir_eq_8_inst0__in1;
  wire  coreir_eq_8_inst0__out;
  coreir_eq #(.width(8)) coreir_eq_8_inst0(
    .in0(coreir_eq_8_inst0__in0),
    .in1(coreir_eq_8_inst0__in1),
    .out(coreir_eq_8_inst0__out)
  );

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__ASYNCRESET = reset;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CE = and_inst0__out;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CLK = clk;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__I[0] = config_data[0];

  assign O[0:0] = Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__O[0:0];

  assign and_inst0__in0 = coreir_eq_8_inst0__out;

  assign and_inst0__in1 = config_en;

  assign coreir_eq_8_inst0__in1[7:0] = const_25_8__out[7:0];

  assign coreir_eq_8_inst0__in0[7:0] = config_addr[7:0];


endmodule  // ConfigRegister_1_8_32_25

module ConfigRegister_1_8_32_23 (
  output [0:0] O,
  input  clk,
  input [7:0] config_addr,
  input [31:0] config_data,
  input  config_en,
  input  reset
);


  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__ASYNCRESET;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CE;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CLK;
  wire [0:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__I;
  wire [0:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__O;
  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1 Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0(
    .ASYNCRESET(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__ASYNCRESET),
    .CE(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CE),
    .CLK(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CLK),
    .I(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__I),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__O)
  );

  wire  and_inst0__in0;
  wire  and_inst0__in1;
  wire  and_inst0__out;
  corebit_and and_inst0(
    .in0(and_inst0__in0),
    .in1(and_inst0__in1),
    .out(and_inst0__out)
  );

  // Instancing generated Module: coreir.const(width:8)
  wire [7:0] const_23_8__out;
  coreir_const #(.value(8'h17),.width(8)) const_23_8(
    .out(const_23_8__out)
  );

  // Instancing generated Module: coreir.eq(width:8)
  wire [7:0] coreir_eq_8_inst0__in0;
  wire [7:0] coreir_eq_8_inst0__in1;
  wire  coreir_eq_8_inst0__out;
  coreir_eq #(.width(8)) coreir_eq_8_inst0(
    .in0(coreir_eq_8_inst0__in0),
    .in1(coreir_eq_8_inst0__in1),
    .out(coreir_eq_8_inst0__out)
  );

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__ASYNCRESET = reset;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CE = and_inst0__out;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CLK = clk;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__I[0] = config_data[0];

  assign O[0:0] = Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__O[0:0];

  assign and_inst0__in0 = coreir_eq_8_inst0__out;

  assign and_inst0__in1 = config_en;

  assign coreir_eq_8_inst0__in1[7:0] = const_23_8__out[7:0];

  assign coreir_eq_8_inst0__in0[7:0] = config_addr[7:0];


endmodule  // ConfigRegister_1_8_32_23

module ConfigRegister_1_8_32_21 (
  output [0:0] O,
  input  clk,
  input [7:0] config_addr,
  input [31:0] config_data,
  input  config_en,
  input  reset
);


  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__ASYNCRESET;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CE;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CLK;
  wire [0:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__I;
  wire [0:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__O;
  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1 Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0(
    .ASYNCRESET(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__ASYNCRESET),
    .CE(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CE),
    .CLK(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CLK),
    .I(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__I),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__O)
  );

  wire  and_inst0__in0;
  wire  and_inst0__in1;
  wire  and_inst0__out;
  corebit_and and_inst0(
    .in0(and_inst0__in0),
    .in1(and_inst0__in1),
    .out(and_inst0__out)
  );

  // Instancing generated Module: coreir.const(width:8)
  wire [7:0] const_21_8__out;
  coreir_const #(.value(8'h15),.width(8)) const_21_8(
    .out(const_21_8__out)
  );

  // Instancing generated Module: coreir.eq(width:8)
  wire [7:0] coreir_eq_8_inst0__in0;
  wire [7:0] coreir_eq_8_inst0__in1;
  wire  coreir_eq_8_inst0__out;
  coreir_eq #(.width(8)) coreir_eq_8_inst0(
    .in0(coreir_eq_8_inst0__in0),
    .in1(coreir_eq_8_inst0__in1),
    .out(coreir_eq_8_inst0__out)
  );

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__ASYNCRESET = reset;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CE = and_inst0__out;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CLK = clk;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__I[0] = config_data[0];

  assign O[0:0] = Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__O[0:0];

  assign and_inst0__in0 = coreir_eq_8_inst0__out;

  assign and_inst0__in1 = config_en;

  assign coreir_eq_8_inst0__in1[7:0] = const_21_8__out[7:0];

  assign coreir_eq_8_inst0__in0[7:0] = config_addr[7:0];


endmodule  // ConfigRegister_1_8_32_21

module ConfigRegister_1_8_32_19 (
  output [0:0] O,
  input  clk,
  input [7:0] config_addr,
  input [31:0] config_data,
  input  config_en,
  input  reset
);


  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__ASYNCRESET;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CE;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CLK;
  wire [0:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__I;
  wire [0:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__O;
  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1 Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0(
    .ASYNCRESET(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__ASYNCRESET),
    .CE(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CE),
    .CLK(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CLK),
    .I(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__I),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__O)
  );

  wire  and_inst0__in0;
  wire  and_inst0__in1;
  wire  and_inst0__out;
  corebit_and and_inst0(
    .in0(and_inst0__in0),
    .in1(and_inst0__in1),
    .out(and_inst0__out)
  );

  // Instancing generated Module: coreir.const(width:8)
  wire [7:0] const_19_8__out;
  coreir_const #(.value(8'h13),.width(8)) const_19_8(
    .out(const_19_8__out)
  );

  // Instancing generated Module: coreir.eq(width:8)
  wire [7:0] coreir_eq_8_inst0__in0;
  wire [7:0] coreir_eq_8_inst0__in1;
  wire  coreir_eq_8_inst0__out;
  coreir_eq #(.width(8)) coreir_eq_8_inst0(
    .in0(coreir_eq_8_inst0__in0),
    .in1(coreir_eq_8_inst0__in1),
    .out(coreir_eq_8_inst0__out)
  );

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__ASYNCRESET = reset;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CE = and_inst0__out;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CLK = clk;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__I[0] = config_data[0];

  assign O[0:0] = Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__O[0:0];

  assign and_inst0__in0 = coreir_eq_8_inst0__out;

  assign and_inst0__in1 = config_en;

  assign coreir_eq_8_inst0__in1[7:0] = const_19_8__out[7:0];

  assign coreir_eq_8_inst0__in0[7:0] = config_addr[7:0];


endmodule  // ConfigRegister_1_8_32_19

module ConfigRegister_1_8_32_17 (
  output [0:0] O,
  input  clk,
  input [7:0] config_addr,
  input [31:0] config_data,
  input  config_en,
  input  reset
);


  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__ASYNCRESET;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CE;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CLK;
  wire [0:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__I;
  wire [0:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__O;
  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1 Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0(
    .ASYNCRESET(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__ASYNCRESET),
    .CE(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CE),
    .CLK(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CLK),
    .I(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__I),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__O)
  );

  wire  and_inst0__in0;
  wire  and_inst0__in1;
  wire  and_inst0__out;
  corebit_and and_inst0(
    .in0(and_inst0__in0),
    .in1(and_inst0__in1),
    .out(and_inst0__out)
  );

  // Instancing generated Module: coreir.const(width:8)
  wire [7:0] const_17_8__out;
  coreir_const #(.value(8'h11),.width(8)) const_17_8(
    .out(const_17_8__out)
  );

  // Instancing generated Module: coreir.eq(width:8)
  wire [7:0] coreir_eq_8_inst0__in0;
  wire [7:0] coreir_eq_8_inst0__in1;
  wire  coreir_eq_8_inst0__out;
  coreir_eq #(.width(8)) coreir_eq_8_inst0(
    .in0(coreir_eq_8_inst0__in0),
    .in1(coreir_eq_8_inst0__in1),
    .out(coreir_eq_8_inst0__out)
  );

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__ASYNCRESET = reset;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CE = and_inst0__out;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CLK = clk;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__I[0] = config_data[0];

  assign O[0:0] = Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__O[0:0];

  assign and_inst0__in0 = coreir_eq_8_inst0__out;

  assign and_inst0__in1 = config_en;

  assign coreir_eq_8_inst0__in1[7:0] = const_17_8__out[7:0];

  assign coreir_eq_8_inst0__in0[7:0] = config_addr[7:0];


endmodule  // ConfigRegister_1_8_32_17

module ConfigRegister_1_8_32_15 (
  output [0:0] O,
  input  clk,
  input [7:0] config_addr,
  input [31:0] config_data,
  input  config_en,
  input  reset
);


  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__ASYNCRESET;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CE;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CLK;
  wire [0:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__I;
  wire [0:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__O;
  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1 Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0(
    .ASYNCRESET(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__ASYNCRESET),
    .CE(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CE),
    .CLK(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CLK),
    .I(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__I),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__O)
  );

  wire  and_inst0__in0;
  wire  and_inst0__in1;
  wire  and_inst0__out;
  corebit_and and_inst0(
    .in0(and_inst0__in0),
    .in1(and_inst0__in1),
    .out(and_inst0__out)
  );

  // Instancing generated Module: coreir.const(width:8)
  wire [7:0] const_15_8__out;
  coreir_const #(.value(8'h0f),.width(8)) const_15_8(
    .out(const_15_8__out)
  );

  // Instancing generated Module: coreir.eq(width:8)
  wire [7:0] coreir_eq_8_inst0__in0;
  wire [7:0] coreir_eq_8_inst0__in1;
  wire  coreir_eq_8_inst0__out;
  coreir_eq #(.width(8)) coreir_eq_8_inst0(
    .in0(coreir_eq_8_inst0__in0),
    .in1(coreir_eq_8_inst0__in1),
    .out(coreir_eq_8_inst0__out)
  );

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__ASYNCRESET = reset;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CE = and_inst0__out;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CLK = clk;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__I[0] = config_data[0];

  assign O[0:0] = Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__O[0:0];

  assign and_inst0__in0 = coreir_eq_8_inst0__out;

  assign and_inst0__in1 = config_en;

  assign coreir_eq_8_inst0__in1[7:0] = const_15_8__out[7:0];

  assign coreir_eq_8_inst0__in0[7:0] = config_addr[7:0];


endmodule  // ConfigRegister_1_8_32_15

module ConfigRegister_1_8_32_13 (
  output [0:0] O,
  input  clk,
  input [7:0] config_addr,
  input [31:0] config_data,
  input  config_en,
  input  reset
);


  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__ASYNCRESET;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CE;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CLK;
  wire [0:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__I;
  wire [0:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__O;
  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1 Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0(
    .ASYNCRESET(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__ASYNCRESET),
    .CE(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CE),
    .CLK(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CLK),
    .I(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__I),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__O)
  );

  wire  and_inst0__in0;
  wire  and_inst0__in1;
  wire  and_inst0__out;
  corebit_and and_inst0(
    .in0(and_inst0__in0),
    .in1(and_inst0__in1),
    .out(and_inst0__out)
  );

  // Instancing generated Module: coreir.const(width:8)
  wire [7:0] const_13_8__out;
  coreir_const #(.value(8'h0d),.width(8)) const_13_8(
    .out(const_13_8__out)
  );

  // Instancing generated Module: coreir.eq(width:8)
  wire [7:0] coreir_eq_8_inst0__in0;
  wire [7:0] coreir_eq_8_inst0__in1;
  wire  coreir_eq_8_inst0__out;
  coreir_eq #(.width(8)) coreir_eq_8_inst0(
    .in0(coreir_eq_8_inst0__in0),
    .in1(coreir_eq_8_inst0__in1),
    .out(coreir_eq_8_inst0__out)
  );

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__ASYNCRESET = reset;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CE = and_inst0__out;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CLK = clk;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__I[0] = config_data[0];

  assign O[0:0] = Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__O[0:0];

  assign and_inst0__in0 = coreir_eq_8_inst0__out;

  assign and_inst0__in1 = config_en;

  assign coreir_eq_8_inst0__in1[7:0] = const_13_8__out[7:0];

  assign coreir_eq_8_inst0__in0[7:0] = config_addr[7:0];


endmodule  // ConfigRegister_1_8_32_13

module ConfigRegister_1_8_32_11 (
  output [0:0] O,
  input  clk,
  input [7:0] config_addr,
  input [31:0] config_data,
  input  config_en,
  input  reset
);


  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__ASYNCRESET;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CE;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CLK;
  wire [0:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__I;
  wire [0:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__O;
  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1 Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0(
    .ASYNCRESET(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__ASYNCRESET),
    .CE(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CE),
    .CLK(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CLK),
    .I(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__I),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__O)
  );

  wire  and_inst0__in0;
  wire  and_inst0__in1;
  wire  and_inst0__out;
  corebit_and and_inst0(
    .in0(and_inst0__in0),
    .in1(and_inst0__in1),
    .out(and_inst0__out)
  );

  // Instancing generated Module: coreir.const(width:8)
  wire [7:0] const_11_8__out;
  coreir_const #(.value(8'h0b),.width(8)) const_11_8(
    .out(const_11_8__out)
  );

  // Instancing generated Module: coreir.eq(width:8)
  wire [7:0] coreir_eq_8_inst0__in0;
  wire [7:0] coreir_eq_8_inst0__in1;
  wire  coreir_eq_8_inst0__out;
  coreir_eq #(.width(8)) coreir_eq_8_inst0(
    .in0(coreir_eq_8_inst0__in0),
    .in1(coreir_eq_8_inst0__in1),
    .out(coreir_eq_8_inst0__out)
  );

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__ASYNCRESET = reset;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CE = and_inst0__out;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CLK = clk;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__I[0] = config_data[0];

  assign O[0:0] = Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__O[0:0];

  assign and_inst0__in0 = coreir_eq_8_inst0__out;

  assign and_inst0__in1 = config_en;

  assign coreir_eq_8_inst0__in1[7:0] = const_11_8__out[7:0];

  assign coreir_eq_8_inst0__in0[7:0] = config_addr[7:0];


endmodule  // ConfigRegister_1_8_32_11

module ConfigRegister_1_8_32_1 (
  output [0:0] O,
  input  clk,
  input [7:0] config_addr,
  input [31:0] config_data,
  input  config_en,
  input  reset
);


  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__ASYNCRESET;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CE;
  wire  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CLK;
  wire [0:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__I;
  wire [0:0] Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__O;
  Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1 Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0(
    .ASYNCRESET(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__ASYNCRESET),
    .CE(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CE),
    .CLK(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CLK),
    .I(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__I),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__O)
  );

  wire  and_inst0__in0;
  wire  and_inst0__in1;
  wire  and_inst0__out;
  corebit_and and_inst0(
    .in0(and_inst0__in0),
    .in1(and_inst0__in1),
    .out(and_inst0__out)
  );

  // Instancing generated Module: coreir.const(width:8)
  wire [7:0] const_1_8__out;
  coreir_const #(.value(8'h01),.width(8)) const_1_8(
    .out(const_1_8__out)
  );

  // Instancing generated Module: coreir.eq(width:8)
  wire [7:0] coreir_eq_8_inst0__in0;
  wire [7:0] coreir_eq_8_inst0__in1;
  wire  coreir_eq_8_inst0__out;
  coreir_eq #(.width(8)) coreir_eq_8_inst0(
    .in0(coreir_eq_8_inst0__in0),
    .in1(coreir_eq_8_inst0__in1),
    .out(coreir_eq_8_inst0__out)
  );

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__ASYNCRESET = reset;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CE = and_inst0__out;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__CLK = clk;

  assign Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__I[0] = config_data[0];

  assign O[0:0] = Register_has_ce_True_has_reset_False_has_async_reset_True_type_Bits_n_1_inst0__O[0:0];

  assign and_inst0__in0 = coreir_eq_8_inst0__out;

  assign and_inst0__in1 = config_en;

  assign coreir_eq_8_inst0__in1[7:0] = const_1_8__out[7:0];

  assign coreir_eq_8_inst0__in0[7:0] = config_addr[7:0];


endmodule  // ConfigRegister_1_8_32_1

module SB_Out_Bits_16___Out_Bits_1__ (
  input  clk,
  input [7:0] config_config_addr,
  input [31:0] config_config_data,
  input [0:0] config_read,
  input [0:0] config_write,
  input [15:0] east_I_layer16_0,
  input [15:0] east_I_layer16_1,
  input [15:0] east_I_layer16_2,
  input [15:0] east_I_layer16_3,
  input [15:0] east_I_layer16_4,
  input [0:0] east_I_layer1_0,
  input [0:0] east_I_layer1_1,
  input [0:0] east_I_layer1_2,
  input [0:0] east_I_layer1_3,
  input [0:0] east_I_layer1_4,
  output [15:0] east_O_layer16_0,
  output [15:0] east_O_layer16_1,
  output [15:0] east_O_layer16_2,
  output [15:0] east_O_layer16_3,
  output [15:0] east_O_layer16_4,
  output [0:0] east_O_layer1_0,
  output [0:0] east_O_layer1_1,
  output [0:0] east_O_layer1_2,
  output [0:0] east_O_layer1_3,
  output [0:0] east_O_layer1_4,
  input [15:0] north_I_layer16_0,
  input [15:0] north_I_layer16_1,
  input [15:0] north_I_layer16_2,
  input [15:0] north_I_layer16_3,
  input [15:0] north_I_layer16_4,
  input [0:0] north_I_layer1_0,
  input [0:0] north_I_layer1_1,
  input [0:0] north_I_layer1_2,
  input [0:0] north_I_layer1_3,
  input [0:0] north_I_layer1_4,
  output [15:0] north_O_layer16_0,
  output [15:0] north_O_layer16_1,
  output [15:0] north_O_layer16_2,
  output [15:0] north_O_layer16_3,
  output [15:0] north_O_layer16_4,
  output [0:0] north_O_layer1_0,
  output [0:0] north_O_layer1_1,
  output [0:0] north_O_layer1_2,
  output [0:0] north_O_layer1_3,
  output [0:0] north_O_layer1_4,
  output [31:0] read_config_data,
  input [15:0] res,
  input [0:0] res_p,
  input  reset,
  input [15:0] south_I_layer16_0,
  input [15:0] south_I_layer16_1,
  input [15:0] south_I_layer16_2,
  input [15:0] south_I_layer16_3,
  input [15:0] south_I_layer16_4,
  input [0:0] south_I_layer1_0,
  input [0:0] south_I_layer1_1,
  input [0:0] south_I_layer1_2,
  input [0:0] south_I_layer1_3,
  input [0:0] south_I_layer1_4,
  output [15:0] south_O_layer16_0,
  output [15:0] south_O_layer16_1,
  output [15:0] south_O_layer16_2,
  output [15:0] south_O_layer16_3,
  output [15:0] south_O_layer16_4,
  output [0:0] south_O_layer1_0,
  output [0:0] south_O_layer1_1,
  output [0:0] south_O_layer1_2,
  output [0:0] south_O_layer1_3,
  output [0:0] south_O_layer1_4,
  input [15:0] west_I_layer16_0,
  input [15:0] west_I_layer16_1,
  input [15:0] west_I_layer16_2,
  input [15:0] west_I_layer16_3,
  input [15:0] west_I_layer16_4,
  input [0:0] west_I_layer1_0,
  input [0:0] west_I_layer1_1,
  input [0:0] west_I_layer1_2,
  input [0:0] west_I_layer1_3,
  input [0:0] west_I_layer1_4,
  output [15:0] west_O_layer16_0,
  output [15:0] west_O_layer16_1,
  output [15:0] west_O_layer16_2,
  output [15:0] west_O_layer16_3,
  output [15:0] west_O_layer16_4,
  output [0:0] west_O_layer1_0,
  output [0:0] west_O_layer1_1,
  output [0:0] west_O_layer1_2,
  output [0:0] west_O_layer1_3,
  output [0:0] west_O_layer1_4
);


  wire [0:0] ConfigRegister_1_8_32_11_inst0__O;
  wire  ConfigRegister_1_8_32_11_inst0__clk;
  wire [7:0] ConfigRegister_1_8_32_11_inst0__config_addr;
  wire [31:0] ConfigRegister_1_8_32_11_inst0__config_data;
  wire  ConfigRegister_1_8_32_11_inst0__config_en;
  wire  ConfigRegister_1_8_32_11_inst0__reset;
  ConfigRegister_1_8_32_11 ConfigRegister_1_8_32_11_inst0(
    .O(ConfigRegister_1_8_32_11_inst0__O),
    .clk(ConfigRegister_1_8_32_11_inst0__clk),
    .config_addr(ConfigRegister_1_8_32_11_inst0__config_addr),
    .config_data(ConfigRegister_1_8_32_11_inst0__config_data),
    .config_en(ConfigRegister_1_8_32_11_inst0__config_en),
    .reset(ConfigRegister_1_8_32_11_inst0__reset)
  );

  wire [0:0] ConfigRegister_1_8_32_13_inst0__O;
  wire  ConfigRegister_1_8_32_13_inst0__clk;
  wire [7:0] ConfigRegister_1_8_32_13_inst0__config_addr;
  wire [31:0] ConfigRegister_1_8_32_13_inst0__config_data;
  wire  ConfigRegister_1_8_32_13_inst0__config_en;
  wire  ConfigRegister_1_8_32_13_inst0__reset;
  ConfigRegister_1_8_32_13 ConfigRegister_1_8_32_13_inst0(
    .O(ConfigRegister_1_8_32_13_inst0__O),
    .clk(ConfigRegister_1_8_32_13_inst0__clk),
    .config_addr(ConfigRegister_1_8_32_13_inst0__config_addr),
    .config_data(ConfigRegister_1_8_32_13_inst0__config_data),
    .config_en(ConfigRegister_1_8_32_13_inst0__config_en),
    .reset(ConfigRegister_1_8_32_13_inst0__reset)
  );

  wire [0:0] ConfigRegister_1_8_32_15_inst0__O;
  wire  ConfigRegister_1_8_32_15_inst0__clk;
  wire [7:0] ConfigRegister_1_8_32_15_inst0__config_addr;
  wire [31:0] ConfigRegister_1_8_32_15_inst0__config_data;
  wire  ConfigRegister_1_8_32_15_inst0__config_en;
  wire  ConfigRegister_1_8_32_15_inst0__reset;
  ConfigRegister_1_8_32_15 ConfigRegister_1_8_32_15_inst0(
    .O(ConfigRegister_1_8_32_15_inst0__O),
    .clk(ConfigRegister_1_8_32_15_inst0__clk),
    .config_addr(ConfigRegister_1_8_32_15_inst0__config_addr),
    .config_data(ConfigRegister_1_8_32_15_inst0__config_data),
    .config_en(ConfigRegister_1_8_32_15_inst0__config_en),
    .reset(ConfigRegister_1_8_32_15_inst0__reset)
  );

  wire [0:0] ConfigRegister_1_8_32_17_inst0__O;
  wire  ConfigRegister_1_8_32_17_inst0__clk;
  wire [7:0] ConfigRegister_1_8_32_17_inst0__config_addr;
  wire [31:0] ConfigRegister_1_8_32_17_inst0__config_data;
  wire  ConfigRegister_1_8_32_17_inst0__config_en;
  wire  ConfigRegister_1_8_32_17_inst0__reset;
  ConfigRegister_1_8_32_17 ConfigRegister_1_8_32_17_inst0(
    .O(ConfigRegister_1_8_32_17_inst0__O),
    .clk(ConfigRegister_1_8_32_17_inst0__clk),
    .config_addr(ConfigRegister_1_8_32_17_inst0__config_addr),
    .config_data(ConfigRegister_1_8_32_17_inst0__config_data),
    .config_en(ConfigRegister_1_8_32_17_inst0__config_en),
    .reset(ConfigRegister_1_8_32_17_inst0__reset)
  );

  wire [0:0] ConfigRegister_1_8_32_19_inst0__O;
  wire  ConfigRegister_1_8_32_19_inst0__clk;
  wire [7:0] ConfigRegister_1_8_32_19_inst0__config_addr;
  wire [31:0] ConfigRegister_1_8_32_19_inst0__config_data;
  wire  ConfigRegister_1_8_32_19_inst0__config_en;
  wire  ConfigRegister_1_8_32_19_inst0__reset;
  ConfigRegister_1_8_32_19 ConfigRegister_1_8_32_19_inst0(
    .O(ConfigRegister_1_8_32_19_inst0__O),
    .clk(ConfigRegister_1_8_32_19_inst0__clk),
    .config_addr(ConfigRegister_1_8_32_19_inst0__config_addr),
    .config_data(ConfigRegister_1_8_32_19_inst0__config_data),
    .config_en(ConfigRegister_1_8_32_19_inst0__config_en),
    .reset(ConfigRegister_1_8_32_19_inst0__reset)
  );

  wire [0:0] ConfigRegister_1_8_32_1_inst0__O;
  wire  ConfigRegister_1_8_32_1_inst0__clk;
  wire [7:0] ConfigRegister_1_8_32_1_inst0__config_addr;
  wire [31:0] ConfigRegister_1_8_32_1_inst0__config_data;
  wire  ConfigRegister_1_8_32_1_inst0__config_en;
  wire  ConfigRegister_1_8_32_1_inst0__reset;
  ConfigRegister_1_8_32_1 ConfigRegister_1_8_32_1_inst0(
    .O(ConfigRegister_1_8_32_1_inst0__O),
    .clk(ConfigRegister_1_8_32_1_inst0__clk),
    .config_addr(ConfigRegister_1_8_32_1_inst0__config_addr),
    .config_data(ConfigRegister_1_8_32_1_inst0__config_data),
    .config_en(ConfigRegister_1_8_32_1_inst0__config_en),
    .reset(ConfigRegister_1_8_32_1_inst0__reset)
  );

  wire [0:0] ConfigRegister_1_8_32_21_inst0__O;
  wire  ConfigRegister_1_8_32_21_inst0__clk;
  wire [7:0] ConfigRegister_1_8_32_21_inst0__config_addr;
  wire [31:0] ConfigRegister_1_8_32_21_inst0__config_data;
  wire  ConfigRegister_1_8_32_21_inst0__config_en;
  wire  ConfigRegister_1_8_32_21_inst0__reset;
  ConfigRegister_1_8_32_21 ConfigRegister_1_8_32_21_inst0(
    .O(ConfigRegister_1_8_32_21_inst0__O),
    .clk(ConfigRegister_1_8_32_21_inst0__clk),
    .config_addr(ConfigRegister_1_8_32_21_inst0__config_addr),
    .config_data(ConfigRegister_1_8_32_21_inst0__config_data),
    .config_en(ConfigRegister_1_8_32_21_inst0__config_en),
    .reset(ConfigRegister_1_8_32_21_inst0__reset)
  );

  wire [0:0] ConfigRegister_1_8_32_23_inst0__O;
  wire  ConfigRegister_1_8_32_23_inst0__clk;
  wire [7:0] ConfigRegister_1_8_32_23_inst0__config_addr;
  wire [31:0] ConfigRegister_1_8_32_23_inst0__config_data;
  wire  ConfigRegister_1_8_32_23_inst0__config_en;
  wire  ConfigRegister_1_8_32_23_inst0__reset;
  ConfigRegister_1_8_32_23 ConfigRegister_1_8_32_23_inst0(
    .O(ConfigRegister_1_8_32_23_inst0__O),
    .clk(ConfigRegister_1_8_32_23_inst0__clk),
    .config_addr(ConfigRegister_1_8_32_23_inst0__config_addr),
    .config_data(ConfigRegister_1_8_32_23_inst0__config_data),
    .config_en(ConfigRegister_1_8_32_23_inst0__config_en),
    .reset(ConfigRegister_1_8_32_23_inst0__reset)
  );

  wire [0:0] ConfigRegister_1_8_32_25_inst0__O;
  wire  ConfigRegister_1_8_32_25_inst0__clk;
  wire [7:0] ConfigRegister_1_8_32_25_inst0__config_addr;
  wire [31:0] ConfigRegister_1_8_32_25_inst0__config_data;
  wire  ConfigRegister_1_8_32_25_inst0__config_en;
  wire  ConfigRegister_1_8_32_25_inst0__reset;
  ConfigRegister_1_8_32_25 ConfigRegister_1_8_32_25_inst0(
    .O(ConfigRegister_1_8_32_25_inst0__O),
    .clk(ConfigRegister_1_8_32_25_inst0__clk),
    .config_addr(ConfigRegister_1_8_32_25_inst0__config_addr),
    .config_data(ConfigRegister_1_8_32_25_inst0__config_data),
    .config_en(ConfigRegister_1_8_32_25_inst0__config_en),
    .reset(ConfigRegister_1_8_32_25_inst0__reset)
  );

  wire [0:0] ConfigRegister_1_8_32_27_inst0__O;
  wire  ConfigRegister_1_8_32_27_inst0__clk;
  wire [7:0] ConfigRegister_1_8_32_27_inst0__config_addr;
  wire [31:0] ConfigRegister_1_8_32_27_inst0__config_data;
  wire  ConfigRegister_1_8_32_27_inst0__config_en;
  wire  ConfigRegister_1_8_32_27_inst0__reset;
  ConfigRegister_1_8_32_27 ConfigRegister_1_8_32_27_inst0(
    .O(ConfigRegister_1_8_32_27_inst0__O),
    .clk(ConfigRegister_1_8_32_27_inst0__clk),
    .config_addr(ConfigRegister_1_8_32_27_inst0__config_addr),
    .config_data(ConfigRegister_1_8_32_27_inst0__config_data),
    .config_en(ConfigRegister_1_8_32_27_inst0__config_en),
    .reset(ConfigRegister_1_8_32_27_inst0__reset)
  );

  wire [0:0] ConfigRegister_1_8_32_29_inst0__O;
  wire  ConfigRegister_1_8_32_29_inst0__clk;
  wire [7:0] ConfigRegister_1_8_32_29_inst0__config_addr;
  wire [31:0] ConfigRegister_1_8_32_29_inst0__config_data;
  wire  ConfigRegister_1_8_32_29_inst0__config_en;
  wire  ConfigRegister_1_8_32_29_inst0__reset;
  ConfigRegister_1_8_32_29 ConfigRegister_1_8_32_29_inst0(
    .O(ConfigRegister_1_8_32_29_inst0__O),
    .clk(ConfigRegister_1_8_32_29_inst0__clk),
    .config_addr(ConfigRegister_1_8_32_29_inst0__config_addr),
    .config_data(ConfigRegister_1_8_32_29_inst0__config_data),
    .config_en(ConfigRegister_1_8_32_29_inst0__config_en),
    .reset(ConfigRegister_1_8_32_29_inst0__reset)
  );

  wire [0:0] ConfigRegister_1_8_32_31_inst0__O;
  wire  ConfigRegister_1_8_32_31_inst0__clk;
  wire [7:0] ConfigRegister_1_8_32_31_inst0__config_addr;
  wire [31:0] ConfigRegister_1_8_32_31_inst0__config_data;
  wire  ConfigRegister_1_8_32_31_inst0__config_en;
  wire  ConfigRegister_1_8_32_31_inst0__reset;
  ConfigRegister_1_8_32_31 ConfigRegister_1_8_32_31_inst0(
    .O(ConfigRegister_1_8_32_31_inst0__O),
    .clk(ConfigRegister_1_8_32_31_inst0__clk),
    .config_addr(ConfigRegister_1_8_32_31_inst0__config_addr),
    .config_data(ConfigRegister_1_8_32_31_inst0__config_data),
    .config_en(ConfigRegister_1_8_32_31_inst0__config_en),
    .reset(ConfigRegister_1_8_32_31_inst0__reset)
  );

  wire [0:0] ConfigRegister_1_8_32_33_inst0__O;
  wire  ConfigRegister_1_8_32_33_inst0__clk;
  wire [7:0] ConfigRegister_1_8_32_33_inst0__config_addr;
  wire [31:0] ConfigRegister_1_8_32_33_inst0__config_data;
  wire  ConfigRegister_1_8_32_33_inst0__config_en;
  wire  ConfigRegister_1_8_32_33_inst0__reset;
  ConfigRegister_1_8_32_33 ConfigRegister_1_8_32_33_inst0(
    .O(ConfigRegister_1_8_32_33_inst0__O),
    .clk(ConfigRegister_1_8_32_33_inst0__clk),
    .config_addr(ConfigRegister_1_8_32_33_inst0__config_addr),
    .config_data(ConfigRegister_1_8_32_33_inst0__config_data),
    .config_en(ConfigRegister_1_8_32_33_inst0__config_en),
    .reset(ConfigRegister_1_8_32_33_inst0__reset)
  );

  wire [0:0] ConfigRegister_1_8_32_35_inst0__O;
  wire  ConfigRegister_1_8_32_35_inst0__clk;
  wire [7:0] ConfigRegister_1_8_32_35_inst0__config_addr;
  wire [31:0] ConfigRegister_1_8_32_35_inst0__config_data;
  wire  ConfigRegister_1_8_32_35_inst0__config_en;
  wire  ConfigRegister_1_8_32_35_inst0__reset;
  ConfigRegister_1_8_32_35 ConfigRegister_1_8_32_35_inst0(
    .O(ConfigRegister_1_8_32_35_inst0__O),
    .clk(ConfigRegister_1_8_32_35_inst0__clk),
    .config_addr(ConfigRegister_1_8_32_35_inst0__config_addr),
    .config_data(ConfigRegister_1_8_32_35_inst0__config_data),
    .config_en(ConfigRegister_1_8_32_35_inst0__config_en),
    .reset(ConfigRegister_1_8_32_35_inst0__reset)
  );

  wire [0:0] ConfigRegister_1_8_32_37_inst0__O;
  wire  ConfigRegister_1_8_32_37_inst0__clk;
  wire [7:0] ConfigRegister_1_8_32_37_inst0__config_addr;
  wire [31:0] ConfigRegister_1_8_32_37_inst0__config_data;
  wire  ConfigRegister_1_8_32_37_inst0__config_en;
  wire  ConfigRegister_1_8_32_37_inst0__reset;
  ConfigRegister_1_8_32_37 ConfigRegister_1_8_32_37_inst0(
    .O(ConfigRegister_1_8_32_37_inst0__O),
    .clk(ConfigRegister_1_8_32_37_inst0__clk),
    .config_addr(ConfigRegister_1_8_32_37_inst0__config_addr),
    .config_data(ConfigRegister_1_8_32_37_inst0__config_data),
    .config_en(ConfigRegister_1_8_32_37_inst0__config_en),
    .reset(ConfigRegister_1_8_32_37_inst0__reset)
  );

  wire [0:0] ConfigRegister_1_8_32_39_inst0__O;
  wire  ConfigRegister_1_8_32_39_inst0__clk;
  wire [7:0] ConfigRegister_1_8_32_39_inst0__config_addr;
  wire [31:0] ConfigRegister_1_8_32_39_inst0__config_data;
  wire  ConfigRegister_1_8_32_39_inst0__config_en;
  wire  ConfigRegister_1_8_32_39_inst0__reset;
  ConfigRegister_1_8_32_39 ConfigRegister_1_8_32_39_inst0(
    .O(ConfigRegister_1_8_32_39_inst0__O),
    .clk(ConfigRegister_1_8_32_39_inst0__clk),
    .config_addr(ConfigRegister_1_8_32_39_inst0__config_addr),
    .config_data(ConfigRegister_1_8_32_39_inst0__config_data),
    .config_en(ConfigRegister_1_8_32_39_inst0__config_en),
    .reset(ConfigRegister_1_8_32_39_inst0__reset)
  );

  wire [0:0] ConfigRegister_1_8_32_3_inst0__O;
  wire  ConfigRegister_1_8_32_3_inst0__clk;
  wire [7:0] ConfigRegister_1_8_32_3_inst0__config_addr;
  wire [31:0] ConfigRegister_1_8_32_3_inst0__config_data;
  wire  ConfigRegister_1_8_32_3_inst0__config_en;
  wire  ConfigRegister_1_8_32_3_inst0__reset;
  ConfigRegister_1_8_32_3 ConfigRegister_1_8_32_3_inst0(
    .O(ConfigRegister_1_8_32_3_inst0__O),
    .clk(ConfigRegister_1_8_32_3_inst0__clk),
    .config_addr(ConfigRegister_1_8_32_3_inst0__config_addr),
    .config_data(ConfigRegister_1_8_32_3_inst0__config_data),
    .config_en(ConfigRegister_1_8_32_3_inst0__config_en),
    .reset(ConfigRegister_1_8_32_3_inst0__reset)
  );

  wire [0:0] ConfigRegister_1_8_32_41_inst0__O;
  wire  ConfigRegister_1_8_32_41_inst0__clk;
  wire [7:0] ConfigRegister_1_8_32_41_inst0__config_addr;
  wire [31:0] ConfigRegister_1_8_32_41_inst0__config_data;
  wire  ConfigRegister_1_8_32_41_inst0__config_en;
  wire  ConfigRegister_1_8_32_41_inst0__reset;
  ConfigRegister_1_8_32_41 ConfigRegister_1_8_32_41_inst0(
    .O(ConfigRegister_1_8_32_41_inst0__O),
    .clk(ConfigRegister_1_8_32_41_inst0__clk),
    .config_addr(ConfigRegister_1_8_32_41_inst0__config_addr),
    .config_data(ConfigRegister_1_8_32_41_inst0__config_data),
    .config_en(ConfigRegister_1_8_32_41_inst0__config_en),
    .reset(ConfigRegister_1_8_32_41_inst0__reset)
  );

  wire [0:0] ConfigRegister_1_8_32_43_inst0__O;
  wire  ConfigRegister_1_8_32_43_inst0__clk;
  wire [7:0] ConfigRegister_1_8_32_43_inst0__config_addr;
  wire [31:0] ConfigRegister_1_8_32_43_inst0__config_data;
  wire  ConfigRegister_1_8_32_43_inst0__config_en;
  wire  ConfigRegister_1_8_32_43_inst0__reset;
  ConfigRegister_1_8_32_43 ConfigRegister_1_8_32_43_inst0(
    .O(ConfigRegister_1_8_32_43_inst0__O),
    .clk(ConfigRegister_1_8_32_43_inst0__clk),
    .config_addr(ConfigRegister_1_8_32_43_inst0__config_addr),
    .config_data(ConfigRegister_1_8_32_43_inst0__config_data),
    .config_en(ConfigRegister_1_8_32_43_inst0__config_en),
    .reset(ConfigRegister_1_8_32_43_inst0__reset)
  );

  wire [0:0] ConfigRegister_1_8_32_45_inst0__O;
  wire  ConfigRegister_1_8_32_45_inst0__clk;
  wire [7:0] ConfigRegister_1_8_32_45_inst0__config_addr;
  wire [31:0] ConfigRegister_1_8_32_45_inst0__config_data;
  wire  ConfigRegister_1_8_32_45_inst0__config_en;
  wire  ConfigRegister_1_8_32_45_inst0__reset;
  ConfigRegister_1_8_32_45 ConfigRegister_1_8_32_45_inst0(
    .O(ConfigRegister_1_8_32_45_inst0__O),
    .clk(ConfigRegister_1_8_32_45_inst0__clk),
    .config_addr(ConfigRegister_1_8_32_45_inst0__config_addr),
    .config_data(ConfigRegister_1_8_32_45_inst0__config_data),
    .config_en(ConfigRegister_1_8_32_45_inst0__config_en),
    .reset(ConfigRegister_1_8_32_45_inst0__reset)
  );

  wire [0:0] ConfigRegister_1_8_32_47_inst0__O;
  wire  ConfigRegister_1_8_32_47_inst0__clk;
  wire [7:0] ConfigRegister_1_8_32_47_inst0__config_addr;
  wire [31:0] ConfigRegister_1_8_32_47_inst0__config_data;
  wire  ConfigRegister_1_8_32_47_inst0__config_en;
  wire  ConfigRegister_1_8_32_47_inst0__reset;
  ConfigRegister_1_8_32_47 ConfigRegister_1_8_32_47_inst0(
    .O(ConfigRegister_1_8_32_47_inst0__O),
    .clk(ConfigRegister_1_8_32_47_inst0__clk),
    .config_addr(ConfigRegister_1_8_32_47_inst0__config_addr),
    .config_data(ConfigRegister_1_8_32_47_inst0__config_data),
    .config_en(ConfigRegister_1_8_32_47_inst0__config_en),
    .reset(ConfigRegister_1_8_32_47_inst0__reset)
  );

  wire [0:0] ConfigRegister_1_8_32_49_inst0__O;
  wire  ConfigRegister_1_8_32_49_inst0__clk;
  wire [7:0] ConfigRegister_1_8_32_49_inst0__config_addr;
  wire [31:0] ConfigRegister_1_8_32_49_inst0__config_data;
  wire  ConfigRegister_1_8_32_49_inst0__config_en;
  wire  ConfigRegister_1_8_32_49_inst0__reset;
  ConfigRegister_1_8_32_49 ConfigRegister_1_8_32_49_inst0(
    .O(ConfigRegister_1_8_32_49_inst0__O),
    .clk(ConfigRegister_1_8_32_49_inst0__clk),
    .config_addr(ConfigRegister_1_8_32_49_inst0__config_addr),
    .config_data(ConfigRegister_1_8_32_49_inst0__config_data),
    .config_en(ConfigRegister_1_8_32_49_inst0__config_en),
    .reset(ConfigRegister_1_8_32_49_inst0__reset)
  );

  wire [0:0] ConfigRegister_1_8_32_51_inst0__O;
  wire  ConfigRegister_1_8_32_51_inst0__clk;
  wire [7:0] ConfigRegister_1_8_32_51_inst0__config_addr;
  wire [31:0] ConfigRegister_1_8_32_51_inst0__config_data;
  wire  ConfigRegister_1_8_32_51_inst0__config_en;
  wire  ConfigRegister_1_8_32_51_inst0__reset;
  ConfigRegister_1_8_32_51 ConfigRegister_1_8_32_51_inst0(
    .O(ConfigRegister_1_8_32_51_inst0__O),
    .clk(ConfigRegister_1_8_32_51_inst0__clk),
    .config_addr(ConfigRegister_1_8_32_51_inst0__config_addr),
    .config_data(ConfigRegister_1_8_32_51_inst0__config_data),
    .config_en(ConfigRegister_1_8_32_51_inst0__config_en),
    .reset(ConfigRegister_1_8_32_51_inst0__reset)
  );

  wire [0:0] ConfigRegister_1_8_32_53_inst0__O;
  wire  ConfigRegister_1_8_32_53_inst0__clk;
  wire [7:0] ConfigRegister_1_8_32_53_inst0__config_addr;
  wire [31:0] ConfigRegister_1_8_32_53_inst0__config_data;
  wire  ConfigRegister_1_8_32_53_inst0__config_en;
  wire  ConfigRegister_1_8_32_53_inst0__reset;
  ConfigRegister_1_8_32_53 ConfigRegister_1_8_32_53_inst0(
    .O(ConfigRegister_1_8_32_53_inst0__O),
    .clk(ConfigRegister_1_8_32_53_inst0__clk),
    .config_addr(ConfigRegister_1_8_32_53_inst0__config_addr),
    .config_data(ConfigRegister_1_8_32_53_inst0__config_data),
    .config_en(ConfigRegister_1_8_32_53_inst0__config_en),
    .reset(ConfigRegister_1_8_32_53_inst0__reset)
  );

  wire [0:0] ConfigRegister_1_8_32_55_inst0__O;
  wire  ConfigRegister_1_8_32_55_inst0__clk;
  wire [7:0] ConfigRegister_1_8_32_55_inst0__config_addr;
  wire [31:0] ConfigRegister_1_8_32_55_inst0__config_data;
  wire  ConfigRegister_1_8_32_55_inst0__config_en;
  wire  ConfigRegister_1_8_32_55_inst0__reset;
  ConfigRegister_1_8_32_55 ConfigRegister_1_8_32_55_inst0(
    .O(ConfigRegister_1_8_32_55_inst0__O),
    .clk(ConfigRegister_1_8_32_55_inst0__clk),
    .config_addr(ConfigRegister_1_8_32_55_inst0__config_addr),
    .config_data(ConfigRegister_1_8_32_55_inst0__config_data),
    .config_en(ConfigRegister_1_8_32_55_inst0__config_en),
    .reset(ConfigRegister_1_8_32_55_inst0__reset)
  );

  wire [0:0] ConfigRegister_1_8_32_57_inst0__O;
  wire  ConfigRegister_1_8_32_57_inst0__clk;
  wire [7:0] ConfigRegister_1_8_32_57_inst0__config_addr;
  wire [31:0] ConfigRegister_1_8_32_57_inst0__config_data;
  wire  ConfigRegister_1_8_32_57_inst0__config_en;
  wire  ConfigRegister_1_8_32_57_inst0__reset;
  ConfigRegister_1_8_32_57 ConfigRegister_1_8_32_57_inst0(
    .O(ConfigRegister_1_8_32_57_inst0__O),
    .clk(ConfigRegister_1_8_32_57_inst0__clk),
    .config_addr(ConfigRegister_1_8_32_57_inst0__config_addr),
    .config_data(ConfigRegister_1_8_32_57_inst0__config_data),
    .config_en(ConfigRegister_1_8_32_57_inst0__config_en),
    .reset(ConfigRegister_1_8_32_57_inst0__reset)
  );

  wire [0:0] ConfigRegister_1_8_32_59_inst0__O;
  wire  ConfigRegister_1_8_32_59_inst0__clk;
  wire [7:0] ConfigRegister_1_8_32_59_inst0__config_addr;
  wire [31:0] ConfigRegister_1_8_32_59_inst0__config_data;
  wire  ConfigRegister_1_8_32_59_inst0__config_en;
  wire  ConfigRegister_1_8_32_59_inst0__reset;
  ConfigRegister_1_8_32_59 ConfigRegister_1_8_32_59_inst0(
    .O(ConfigRegister_1_8_32_59_inst0__O),
    .clk(ConfigRegister_1_8_32_59_inst0__clk),
    .config_addr(ConfigRegister_1_8_32_59_inst0__config_addr),
    .config_data(ConfigRegister_1_8_32_59_inst0__config_data),
    .config_en(ConfigRegister_1_8_32_59_inst0__config_en),
    .reset(ConfigRegister_1_8_32_59_inst0__reset)
  );

  wire [0:0] ConfigRegister_1_8_32_5_inst0__O;
  wire  ConfigRegister_1_8_32_5_inst0__clk;
  wire [7:0] ConfigRegister_1_8_32_5_inst0__config_addr;
  wire [31:0] ConfigRegister_1_8_32_5_inst0__config_data;
  wire  ConfigRegister_1_8_32_5_inst0__config_en;
  wire  ConfigRegister_1_8_32_5_inst0__reset;
  ConfigRegister_1_8_32_5 ConfigRegister_1_8_32_5_inst0(
    .O(ConfigRegister_1_8_32_5_inst0__O),
    .clk(ConfigRegister_1_8_32_5_inst0__clk),
    .config_addr(ConfigRegister_1_8_32_5_inst0__config_addr),
    .config_data(ConfigRegister_1_8_32_5_inst0__config_data),
    .config_en(ConfigRegister_1_8_32_5_inst0__config_en),
    .reset(ConfigRegister_1_8_32_5_inst0__reset)
  );

  wire [0:0] ConfigRegister_1_8_32_61_inst0__O;
  wire  ConfigRegister_1_8_32_61_inst0__clk;
  wire [7:0] ConfigRegister_1_8_32_61_inst0__config_addr;
  wire [31:0] ConfigRegister_1_8_32_61_inst0__config_data;
  wire  ConfigRegister_1_8_32_61_inst0__config_en;
  wire  ConfigRegister_1_8_32_61_inst0__reset;
  ConfigRegister_1_8_32_61 ConfigRegister_1_8_32_61_inst0(
    .O(ConfigRegister_1_8_32_61_inst0__O),
    .clk(ConfigRegister_1_8_32_61_inst0__clk),
    .config_addr(ConfigRegister_1_8_32_61_inst0__config_addr),
    .config_data(ConfigRegister_1_8_32_61_inst0__config_data),
    .config_en(ConfigRegister_1_8_32_61_inst0__config_en),
    .reset(ConfigRegister_1_8_32_61_inst0__reset)
  );

  wire [0:0] ConfigRegister_1_8_32_63_inst0__O;
  wire  ConfigRegister_1_8_32_63_inst0__clk;
  wire [7:0] ConfigRegister_1_8_32_63_inst0__config_addr;
  wire [31:0] ConfigRegister_1_8_32_63_inst0__config_data;
  wire  ConfigRegister_1_8_32_63_inst0__config_en;
  wire  ConfigRegister_1_8_32_63_inst0__reset;
  ConfigRegister_1_8_32_63 ConfigRegister_1_8_32_63_inst0(
    .O(ConfigRegister_1_8_32_63_inst0__O),
    .clk(ConfigRegister_1_8_32_63_inst0__clk),
    .config_addr(ConfigRegister_1_8_32_63_inst0__config_addr),
    .config_data(ConfigRegister_1_8_32_63_inst0__config_data),
    .config_en(ConfigRegister_1_8_32_63_inst0__config_en),
    .reset(ConfigRegister_1_8_32_63_inst0__reset)
  );

  wire [0:0] ConfigRegister_1_8_32_65_inst0__O;
  wire  ConfigRegister_1_8_32_65_inst0__clk;
  wire [7:0] ConfigRegister_1_8_32_65_inst0__config_addr;
  wire [31:0] ConfigRegister_1_8_32_65_inst0__config_data;
  wire  ConfigRegister_1_8_32_65_inst0__config_en;
  wire  ConfigRegister_1_8_32_65_inst0__reset;
  ConfigRegister_1_8_32_65 ConfigRegister_1_8_32_65_inst0(
    .O(ConfigRegister_1_8_32_65_inst0__O),
    .clk(ConfigRegister_1_8_32_65_inst0__clk),
    .config_addr(ConfigRegister_1_8_32_65_inst0__config_addr),
    .config_data(ConfigRegister_1_8_32_65_inst0__config_data),
    .config_en(ConfigRegister_1_8_32_65_inst0__config_en),
    .reset(ConfigRegister_1_8_32_65_inst0__reset)
  );

  wire [0:0] ConfigRegister_1_8_32_67_inst0__O;
  wire  ConfigRegister_1_8_32_67_inst0__clk;
  wire [7:0] ConfigRegister_1_8_32_67_inst0__config_addr;
  wire [31:0] ConfigRegister_1_8_32_67_inst0__config_data;
  wire  ConfigRegister_1_8_32_67_inst0__config_en;
  wire  ConfigRegister_1_8_32_67_inst0__reset;
  ConfigRegister_1_8_32_67 ConfigRegister_1_8_32_67_inst0(
    .O(ConfigRegister_1_8_32_67_inst0__O),
    .clk(ConfigRegister_1_8_32_67_inst0__clk),
    .config_addr(ConfigRegister_1_8_32_67_inst0__config_addr),
    .config_data(ConfigRegister_1_8_32_67_inst0__config_data),
    .config_en(ConfigRegister_1_8_32_67_inst0__config_en),
    .reset(ConfigRegister_1_8_32_67_inst0__reset)
  );

  wire [0:0] ConfigRegister_1_8_32_69_inst0__O;
  wire  ConfigRegister_1_8_32_69_inst0__clk;
  wire [7:0] ConfigRegister_1_8_32_69_inst0__config_addr;
  wire [31:0] ConfigRegister_1_8_32_69_inst0__config_data;
  wire  ConfigRegister_1_8_32_69_inst0__config_en;
  wire  ConfigRegister_1_8_32_69_inst0__reset;
  ConfigRegister_1_8_32_69 ConfigRegister_1_8_32_69_inst0(
    .O(ConfigRegister_1_8_32_69_inst0__O),
    .clk(ConfigRegister_1_8_32_69_inst0__clk),
    .config_addr(ConfigRegister_1_8_32_69_inst0__config_addr),
    .config_data(ConfigRegister_1_8_32_69_inst0__config_data),
    .config_en(ConfigRegister_1_8_32_69_inst0__config_en),
    .reset(ConfigRegister_1_8_32_69_inst0__reset)
  );

  wire [0:0] ConfigRegister_1_8_32_71_inst0__O;
  wire  ConfigRegister_1_8_32_71_inst0__clk;
  wire [7:0] ConfigRegister_1_8_32_71_inst0__config_addr;
  wire [31:0] ConfigRegister_1_8_32_71_inst0__config_data;
  wire  ConfigRegister_1_8_32_71_inst0__config_en;
  wire  ConfigRegister_1_8_32_71_inst0__reset;
  ConfigRegister_1_8_32_71 ConfigRegister_1_8_32_71_inst0(
    .O(ConfigRegister_1_8_32_71_inst0__O),
    .clk(ConfigRegister_1_8_32_71_inst0__clk),
    .config_addr(ConfigRegister_1_8_32_71_inst0__config_addr),
    .config_data(ConfigRegister_1_8_32_71_inst0__config_data),
    .config_en(ConfigRegister_1_8_32_71_inst0__config_en),
    .reset(ConfigRegister_1_8_32_71_inst0__reset)
  );

  wire [0:0] ConfigRegister_1_8_32_73_inst0__O;
  wire  ConfigRegister_1_8_32_73_inst0__clk;
  wire [7:0] ConfigRegister_1_8_32_73_inst0__config_addr;
  wire [31:0] ConfigRegister_1_8_32_73_inst0__config_data;
  wire  ConfigRegister_1_8_32_73_inst0__config_en;
  wire  ConfigRegister_1_8_32_73_inst0__reset;
  ConfigRegister_1_8_32_73 ConfigRegister_1_8_32_73_inst0(
    .O(ConfigRegister_1_8_32_73_inst0__O),
    .clk(ConfigRegister_1_8_32_73_inst0__clk),
    .config_addr(ConfigRegister_1_8_32_73_inst0__config_addr),
    .config_data(ConfigRegister_1_8_32_73_inst0__config_data),
    .config_en(ConfigRegister_1_8_32_73_inst0__config_en),
    .reset(ConfigRegister_1_8_32_73_inst0__reset)
  );

  wire [0:0] ConfigRegister_1_8_32_75_inst0__O;
  wire  ConfigRegister_1_8_32_75_inst0__clk;
  wire [7:0] ConfigRegister_1_8_32_75_inst0__config_addr;
  wire [31:0] ConfigRegister_1_8_32_75_inst0__config_data;
  wire  ConfigRegister_1_8_32_75_inst0__config_en;
  wire  ConfigRegister_1_8_32_75_inst0__reset;
  ConfigRegister_1_8_32_75 ConfigRegister_1_8_32_75_inst0(
    .O(ConfigRegister_1_8_32_75_inst0__O),
    .clk(ConfigRegister_1_8_32_75_inst0__clk),
    .config_addr(ConfigRegister_1_8_32_75_inst0__config_addr),
    .config_data(ConfigRegister_1_8_32_75_inst0__config_data),
    .config_en(ConfigRegister_1_8_32_75_inst0__config_en),
    .reset(ConfigRegister_1_8_32_75_inst0__reset)
  );

  wire [0:0] ConfigRegister_1_8_32_77_inst0__O;
  wire  ConfigRegister_1_8_32_77_inst0__clk;
  wire [7:0] ConfigRegister_1_8_32_77_inst0__config_addr;
  wire [31:0] ConfigRegister_1_8_32_77_inst0__config_data;
  wire  ConfigRegister_1_8_32_77_inst0__config_en;
  wire  ConfigRegister_1_8_32_77_inst0__reset;
  ConfigRegister_1_8_32_77 ConfigRegister_1_8_32_77_inst0(
    .O(ConfigRegister_1_8_32_77_inst0__O),
    .clk(ConfigRegister_1_8_32_77_inst0__clk),
    .config_addr(ConfigRegister_1_8_32_77_inst0__config_addr),
    .config_data(ConfigRegister_1_8_32_77_inst0__config_data),
    .config_en(ConfigRegister_1_8_32_77_inst0__config_en),
    .reset(ConfigRegister_1_8_32_77_inst0__reset)
  );

  wire [0:0] ConfigRegister_1_8_32_79_inst0__O;
  wire  ConfigRegister_1_8_32_79_inst0__clk;
  wire [7:0] ConfigRegister_1_8_32_79_inst0__config_addr;
  wire [31:0] ConfigRegister_1_8_32_79_inst0__config_data;
  wire  ConfigRegister_1_8_32_79_inst0__config_en;
  wire  ConfigRegister_1_8_32_79_inst0__reset;
  ConfigRegister_1_8_32_79 ConfigRegister_1_8_32_79_inst0(
    .O(ConfigRegister_1_8_32_79_inst0__O),
    .clk(ConfigRegister_1_8_32_79_inst0__clk),
    .config_addr(ConfigRegister_1_8_32_79_inst0__config_addr),
    .config_data(ConfigRegister_1_8_32_79_inst0__config_data),
    .config_en(ConfigRegister_1_8_32_79_inst0__config_en),
    .reset(ConfigRegister_1_8_32_79_inst0__reset)
  );

  wire [0:0] ConfigRegister_1_8_32_7_inst0__O;
  wire  ConfigRegister_1_8_32_7_inst0__clk;
  wire [7:0] ConfigRegister_1_8_32_7_inst0__config_addr;
  wire [31:0] ConfigRegister_1_8_32_7_inst0__config_data;
  wire  ConfigRegister_1_8_32_7_inst0__config_en;
  wire  ConfigRegister_1_8_32_7_inst0__reset;
  ConfigRegister_1_8_32_7 ConfigRegister_1_8_32_7_inst0(
    .O(ConfigRegister_1_8_32_7_inst0__O),
    .clk(ConfigRegister_1_8_32_7_inst0__clk),
    .config_addr(ConfigRegister_1_8_32_7_inst0__config_addr),
    .config_data(ConfigRegister_1_8_32_7_inst0__config_data),
    .config_en(ConfigRegister_1_8_32_7_inst0__config_en),
    .reset(ConfigRegister_1_8_32_7_inst0__reset)
  );

  wire [0:0] ConfigRegister_1_8_32_9_inst0__O;
  wire  ConfigRegister_1_8_32_9_inst0__clk;
  wire [7:0] ConfigRegister_1_8_32_9_inst0__config_addr;
  wire [31:0] ConfigRegister_1_8_32_9_inst0__config_data;
  wire  ConfigRegister_1_8_32_9_inst0__config_en;
  wire  ConfigRegister_1_8_32_9_inst0__reset;
  ConfigRegister_1_8_32_9 ConfigRegister_1_8_32_9_inst0(
    .O(ConfigRegister_1_8_32_9_inst0__O),
    .clk(ConfigRegister_1_8_32_9_inst0__clk),
    .config_addr(ConfigRegister_1_8_32_9_inst0__config_addr),
    .config_data(ConfigRegister_1_8_32_9_inst0__config_data),
    .config_en(ConfigRegister_1_8_32_9_inst0__config_en),
    .reset(ConfigRegister_1_8_32_9_inst0__reset)
  );

  wire [1:0] ConfigRegister_2_8_32_0_inst0__O;
  wire  ConfigRegister_2_8_32_0_inst0__clk;
  wire [7:0] ConfigRegister_2_8_32_0_inst0__config_addr;
  wire [31:0] ConfigRegister_2_8_32_0_inst0__config_data;
  wire  ConfigRegister_2_8_32_0_inst0__config_en;
  wire  ConfigRegister_2_8_32_0_inst0__reset;
  ConfigRegister_2_8_32_0 ConfigRegister_2_8_32_0_inst0(
    .O(ConfigRegister_2_8_32_0_inst0__O),
    .clk(ConfigRegister_2_8_32_0_inst0__clk),
    .config_addr(ConfigRegister_2_8_32_0_inst0__config_addr),
    .config_data(ConfigRegister_2_8_32_0_inst0__config_data),
    .config_en(ConfigRegister_2_8_32_0_inst0__config_en),
    .reset(ConfigRegister_2_8_32_0_inst0__reset)
  );

  wire [1:0] ConfigRegister_2_8_32_10_inst0__O;
  wire  ConfigRegister_2_8_32_10_inst0__clk;
  wire [7:0] ConfigRegister_2_8_32_10_inst0__config_addr;
  wire [31:0] ConfigRegister_2_8_32_10_inst0__config_data;
  wire  ConfigRegister_2_8_32_10_inst0__config_en;
  wire  ConfigRegister_2_8_32_10_inst0__reset;
  ConfigRegister_2_8_32_10 ConfigRegister_2_8_32_10_inst0(
    .O(ConfigRegister_2_8_32_10_inst0__O),
    .clk(ConfigRegister_2_8_32_10_inst0__clk),
    .config_addr(ConfigRegister_2_8_32_10_inst0__config_addr),
    .config_data(ConfigRegister_2_8_32_10_inst0__config_data),
    .config_en(ConfigRegister_2_8_32_10_inst0__config_en),
    .reset(ConfigRegister_2_8_32_10_inst0__reset)
  );

  wire [1:0] ConfigRegister_2_8_32_12_inst0__O;
  wire  ConfigRegister_2_8_32_12_inst0__clk;
  wire [7:0] ConfigRegister_2_8_32_12_inst0__config_addr;
  wire [31:0] ConfigRegister_2_8_32_12_inst0__config_data;
  wire  ConfigRegister_2_8_32_12_inst0__config_en;
  wire  ConfigRegister_2_8_32_12_inst0__reset;
  ConfigRegister_2_8_32_12 ConfigRegister_2_8_32_12_inst0(
    .O(ConfigRegister_2_8_32_12_inst0__O),
    .clk(ConfigRegister_2_8_32_12_inst0__clk),
    .config_addr(ConfigRegister_2_8_32_12_inst0__config_addr),
    .config_data(ConfigRegister_2_8_32_12_inst0__config_data),
    .config_en(ConfigRegister_2_8_32_12_inst0__config_en),
    .reset(ConfigRegister_2_8_32_12_inst0__reset)
  );

  wire [1:0] ConfigRegister_2_8_32_14_inst0__O;
  wire  ConfigRegister_2_8_32_14_inst0__clk;
  wire [7:0] ConfigRegister_2_8_32_14_inst0__config_addr;
  wire [31:0] ConfigRegister_2_8_32_14_inst0__config_data;
  wire  ConfigRegister_2_8_32_14_inst0__config_en;
  wire  ConfigRegister_2_8_32_14_inst0__reset;
  ConfigRegister_2_8_32_14 ConfigRegister_2_8_32_14_inst0(
    .O(ConfigRegister_2_8_32_14_inst0__O),
    .clk(ConfigRegister_2_8_32_14_inst0__clk),
    .config_addr(ConfigRegister_2_8_32_14_inst0__config_addr),
    .config_data(ConfigRegister_2_8_32_14_inst0__config_data),
    .config_en(ConfigRegister_2_8_32_14_inst0__config_en),
    .reset(ConfigRegister_2_8_32_14_inst0__reset)
  );

  wire [1:0] ConfigRegister_2_8_32_16_inst0__O;
  wire  ConfigRegister_2_8_32_16_inst0__clk;
  wire [7:0] ConfigRegister_2_8_32_16_inst0__config_addr;
  wire [31:0] ConfigRegister_2_8_32_16_inst0__config_data;
  wire  ConfigRegister_2_8_32_16_inst0__config_en;
  wire  ConfigRegister_2_8_32_16_inst0__reset;
  ConfigRegister_2_8_32_16 ConfigRegister_2_8_32_16_inst0(
    .O(ConfigRegister_2_8_32_16_inst0__O),
    .clk(ConfigRegister_2_8_32_16_inst0__clk),
    .config_addr(ConfigRegister_2_8_32_16_inst0__config_addr),
    .config_data(ConfigRegister_2_8_32_16_inst0__config_data),
    .config_en(ConfigRegister_2_8_32_16_inst0__config_en),
    .reset(ConfigRegister_2_8_32_16_inst0__reset)
  );

  wire [1:0] ConfigRegister_2_8_32_18_inst0__O;
  wire  ConfigRegister_2_8_32_18_inst0__clk;
  wire [7:0] ConfigRegister_2_8_32_18_inst0__config_addr;
  wire [31:0] ConfigRegister_2_8_32_18_inst0__config_data;
  wire  ConfigRegister_2_8_32_18_inst0__config_en;
  wire  ConfigRegister_2_8_32_18_inst0__reset;
  ConfigRegister_2_8_32_18 ConfigRegister_2_8_32_18_inst0(
    .O(ConfigRegister_2_8_32_18_inst0__O),
    .clk(ConfigRegister_2_8_32_18_inst0__clk),
    .config_addr(ConfigRegister_2_8_32_18_inst0__config_addr),
    .config_data(ConfigRegister_2_8_32_18_inst0__config_data),
    .config_en(ConfigRegister_2_8_32_18_inst0__config_en),
    .reset(ConfigRegister_2_8_32_18_inst0__reset)
  );

  wire [1:0] ConfigRegister_2_8_32_20_inst0__O;
  wire  ConfigRegister_2_8_32_20_inst0__clk;
  wire [7:0] ConfigRegister_2_8_32_20_inst0__config_addr;
  wire [31:0] ConfigRegister_2_8_32_20_inst0__config_data;
  wire  ConfigRegister_2_8_32_20_inst0__config_en;
  wire  ConfigRegister_2_8_32_20_inst0__reset;
  ConfigRegister_2_8_32_20 ConfigRegister_2_8_32_20_inst0(
    .O(ConfigRegister_2_8_32_20_inst0__O),
    .clk(ConfigRegister_2_8_32_20_inst0__clk),
    .config_addr(ConfigRegister_2_8_32_20_inst0__config_addr),
    .config_data(ConfigRegister_2_8_32_20_inst0__config_data),
    .config_en(ConfigRegister_2_8_32_20_inst0__config_en),
    .reset(ConfigRegister_2_8_32_20_inst0__reset)
  );

  wire [1:0] ConfigRegister_2_8_32_22_inst0__O;
  wire  ConfigRegister_2_8_32_22_inst0__clk;
  wire [7:0] ConfigRegister_2_8_32_22_inst0__config_addr;
  wire [31:0] ConfigRegister_2_8_32_22_inst0__config_data;
  wire  ConfigRegister_2_8_32_22_inst0__config_en;
  wire  ConfigRegister_2_8_32_22_inst0__reset;
  ConfigRegister_2_8_32_22 ConfigRegister_2_8_32_22_inst0(
    .O(ConfigRegister_2_8_32_22_inst0__O),
    .clk(ConfigRegister_2_8_32_22_inst0__clk),
    .config_addr(ConfigRegister_2_8_32_22_inst0__config_addr),
    .config_data(ConfigRegister_2_8_32_22_inst0__config_data),
    .config_en(ConfigRegister_2_8_32_22_inst0__config_en),
    .reset(ConfigRegister_2_8_32_22_inst0__reset)
  );

  wire [1:0] ConfigRegister_2_8_32_24_inst0__O;
  wire  ConfigRegister_2_8_32_24_inst0__clk;
  wire [7:0] ConfigRegister_2_8_32_24_inst0__config_addr;
  wire [31:0] ConfigRegister_2_8_32_24_inst0__config_data;
  wire  ConfigRegister_2_8_32_24_inst0__config_en;
  wire  ConfigRegister_2_8_32_24_inst0__reset;
  ConfigRegister_2_8_32_24 ConfigRegister_2_8_32_24_inst0(
    .O(ConfigRegister_2_8_32_24_inst0__O),
    .clk(ConfigRegister_2_8_32_24_inst0__clk),
    .config_addr(ConfigRegister_2_8_32_24_inst0__config_addr),
    .config_data(ConfigRegister_2_8_32_24_inst0__config_data),
    .config_en(ConfigRegister_2_8_32_24_inst0__config_en),
    .reset(ConfigRegister_2_8_32_24_inst0__reset)
  );

  wire [1:0] ConfigRegister_2_8_32_26_inst0__O;
  wire  ConfigRegister_2_8_32_26_inst0__clk;
  wire [7:0] ConfigRegister_2_8_32_26_inst0__config_addr;
  wire [31:0] ConfigRegister_2_8_32_26_inst0__config_data;
  wire  ConfigRegister_2_8_32_26_inst0__config_en;
  wire  ConfigRegister_2_8_32_26_inst0__reset;
  ConfigRegister_2_8_32_26 ConfigRegister_2_8_32_26_inst0(
    .O(ConfigRegister_2_8_32_26_inst0__O),
    .clk(ConfigRegister_2_8_32_26_inst0__clk),
    .config_addr(ConfigRegister_2_8_32_26_inst0__config_addr),
    .config_data(ConfigRegister_2_8_32_26_inst0__config_data),
    .config_en(ConfigRegister_2_8_32_26_inst0__config_en),
    .reset(ConfigRegister_2_8_32_26_inst0__reset)
  );

  wire [1:0] ConfigRegister_2_8_32_28_inst0__O;
  wire  ConfigRegister_2_8_32_28_inst0__clk;
  wire [7:0] ConfigRegister_2_8_32_28_inst0__config_addr;
  wire [31:0] ConfigRegister_2_8_32_28_inst0__config_data;
  wire  ConfigRegister_2_8_32_28_inst0__config_en;
  wire  ConfigRegister_2_8_32_28_inst0__reset;
  ConfigRegister_2_8_32_28 ConfigRegister_2_8_32_28_inst0(
    .O(ConfigRegister_2_8_32_28_inst0__O),
    .clk(ConfigRegister_2_8_32_28_inst0__clk),
    .config_addr(ConfigRegister_2_8_32_28_inst0__config_addr),
    .config_data(ConfigRegister_2_8_32_28_inst0__config_data),
    .config_en(ConfigRegister_2_8_32_28_inst0__config_en),
    .reset(ConfigRegister_2_8_32_28_inst0__reset)
  );

  wire [1:0] ConfigRegister_2_8_32_2_inst0__O;
  wire  ConfigRegister_2_8_32_2_inst0__clk;
  wire [7:0] ConfigRegister_2_8_32_2_inst0__config_addr;
  wire [31:0] ConfigRegister_2_8_32_2_inst0__config_data;
  wire  ConfigRegister_2_8_32_2_inst0__config_en;
  wire  ConfigRegister_2_8_32_2_inst0__reset;
  ConfigRegister_2_8_32_2 ConfigRegister_2_8_32_2_inst0(
    .O(ConfigRegister_2_8_32_2_inst0__O),
    .clk(ConfigRegister_2_8_32_2_inst0__clk),
    .config_addr(ConfigRegister_2_8_32_2_inst0__config_addr),
    .config_data(ConfigRegister_2_8_32_2_inst0__config_data),
    .config_en(ConfigRegister_2_8_32_2_inst0__config_en),
    .reset(ConfigRegister_2_8_32_2_inst0__reset)
  );

  wire [1:0] ConfigRegister_2_8_32_30_inst0__O;
  wire  ConfigRegister_2_8_32_30_inst0__clk;
  wire [7:0] ConfigRegister_2_8_32_30_inst0__config_addr;
  wire [31:0] ConfigRegister_2_8_32_30_inst0__config_data;
  wire  ConfigRegister_2_8_32_30_inst0__config_en;
  wire  ConfigRegister_2_8_32_30_inst0__reset;
  ConfigRegister_2_8_32_30 ConfigRegister_2_8_32_30_inst0(
    .O(ConfigRegister_2_8_32_30_inst0__O),
    .clk(ConfigRegister_2_8_32_30_inst0__clk),
    .config_addr(ConfigRegister_2_8_32_30_inst0__config_addr),
    .config_data(ConfigRegister_2_8_32_30_inst0__config_data),
    .config_en(ConfigRegister_2_8_32_30_inst0__config_en),
    .reset(ConfigRegister_2_8_32_30_inst0__reset)
  );

  wire [1:0] ConfigRegister_2_8_32_32_inst0__O;
  wire  ConfigRegister_2_8_32_32_inst0__clk;
  wire [7:0] ConfigRegister_2_8_32_32_inst0__config_addr;
  wire [31:0] ConfigRegister_2_8_32_32_inst0__config_data;
  wire  ConfigRegister_2_8_32_32_inst0__config_en;
  wire  ConfigRegister_2_8_32_32_inst0__reset;
  ConfigRegister_2_8_32_32 ConfigRegister_2_8_32_32_inst0(
    .O(ConfigRegister_2_8_32_32_inst0__O),
    .clk(ConfigRegister_2_8_32_32_inst0__clk),
    .config_addr(ConfigRegister_2_8_32_32_inst0__config_addr),
    .config_data(ConfigRegister_2_8_32_32_inst0__config_data),
    .config_en(ConfigRegister_2_8_32_32_inst0__config_en),
    .reset(ConfigRegister_2_8_32_32_inst0__reset)
  );

  wire [1:0] ConfigRegister_2_8_32_34_inst0__O;
  wire  ConfigRegister_2_8_32_34_inst0__clk;
  wire [7:0] ConfigRegister_2_8_32_34_inst0__config_addr;
  wire [31:0] ConfigRegister_2_8_32_34_inst0__config_data;
  wire  ConfigRegister_2_8_32_34_inst0__config_en;
  wire  ConfigRegister_2_8_32_34_inst0__reset;
  ConfigRegister_2_8_32_34 ConfigRegister_2_8_32_34_inst0(
    .O(ConfigRegister_2_8_32_34_inst0__O),
    .clk(ConfigRegister_2_8_32_34_inst0__clk),
    .config_addr(ConfigRegister_2_8_32_34_inst0__config_addr),
    .config_data(ConfigRegister_2_8_32_34_inst0__config_data),
    .config_en(ConfigRegister_2_8_32_34_inst0__config_en),
    .reset(ConfigRegister_2_8_32_34_inst0__reset)
  );

  wire [1:0] ConfigRegister_2_8_32_36_inst0__O;
  wire  ConfigRegister_2_8_32_36_inst0__clk;
  wire [7:0] ConfigRegister_2_8_32_36_inst0__config_addr;
  wire [31:0] ConfigRegister_2_8_32_36_inst0__config_data;
  wire  ConfigRegister_2_8_32_36_inst0__config_en;
  wire  ConfigRegister_2_8_32_36_inst0__reset;
  ConfigRegister_2_8_32_36 ConfigRegister_2_8_32_36_inst0(
    .O(ConfigRegister_2_8_32_36_inst0__O),
    .clk(ConfigRegister_2_8_32_36_inst0__clk),
    .config_addr(ConfigRegister_2_8_32_36_inst0__config_addr),
    .config_data(ConfigRegister_2_8_32_36_inst0__config_data),
    .config_en(ConfigRegister_2_8_32_36_inst0__config_en),
    .reset(ConfigRegister_2_8_32_36_inst0__reset)
  );

  wire [1:0] ConfigRegister_2_8_32_38_inst0__O;
  wire  ConfigRegister_2_8_32_38_inst0__clk;
  wire [7:0] ConfigRegister_2_8_32_38_inst0__config_addr;
  wire [31:0] ConfigRegister_2_8_32_38_inst0__config_data;
  wire  ConfigRegister_2_8_32_38_inst0__config_en;
  wire  ConfigRegister_2_8_32_38_inst0__reset;
  ConfigRegister_2_8_32_38 ConfigRegister_2_8_32_38_inst0(
    .O(ConfigRegister_2_8_32_38_inst0__O),
    .clk(ConfigRegister_2_8_32_38_inst0__clk),
    .config_addr(ConfigRegister_2_8_32_38_inst0__config_addr),
    .config_data(ConfigRegister_2_8_32_38_inst0__config_data),
    .config_en(ConfigRegister_2_8_32_38_inst0__config_en),
    .reset(ConfigRegister_2_8_32_38_inst0__reset)
  );

  wire [1:0] ConfigRegister_2_8_32_40_inst0__O;
  wire  ConfigRegister_2_8_32_40_inst0__clk;
  wire [7:0] ConfigRegister_2_8_32_40_inst0__config_addr;
  wire [31:0] ConfigRegister_2_8_32_40_inst0__config_data;
  wire  ConfigRegister_2_8_32_40_inst0__config_en;
  wire  ConfigRegister_2_8_32_40_inst0__reset;
  ConfigRegister_2_8_32_40 ConfigRegister_2_8_32_40_inst0(
    .O(ConfigRegister_2_8_32_40_inst0__O),
    .clk(ConfigRegister_2_8_32_40_inst0__clk),
    .config_addr(ConfigRegister_2_8_32_40_inst0__config_addr),
    .config_data(ConfigRegister_2_8_32_40_inst0__config_data),
    .config_en(ConfigRegister_2_8_32_40_inst0__config_en),
    .reset(ConfigRegister_2_8_32_40_inst0__reset)
  );

  wire [1:0] ConfigRegister_2_8_32_42_inst0__O;
  wire  ConfigRegister_2_8_32_42_inst0__clk;
  wire [7:0] ConfigRegister_2_8_32_42_inst0__config_addr;
  wire [31:0] ConfigRegister_2_8_32_42_inst0__config_data;
  wire  ConfigRegister_2_8_32_42_inst0__config_en;
  wire  ConfigRegister_2_8_32_42_inst0__reset;
  ConfigRegister_2_8_32_42 ConfigRegister_2_8_32_42_inst0(
    .O(ConfigRegister_2_8_32_42_inst0__O),
    .clk(ConfigRegister_2_8_32_42_inst0__clk),
    .config_addr(ConfigRegister_2_8_32_42_inst0__config_addr),
    .config_data(ConfigRegister_2_8_32_42_inst0__config_data),
    .config_en(ConfigRegister_2_8_32_42_inst0__config_en),
    .reset(ConfigRegister_2_8_32_42_inst0__reset)
  );

  wire [1:0] ConfigRegister_2_8_32_44_inst0__O;
  wire  ConfigRegister_2_8_32_44_inst0__clk;
  wire [7:0] ConfigRegister_2_8_32_44_inst0__config_addr;
  wire [31:0] ConfigRegister_2_8_32_44_inst0__config_data;
  wire  ConfigRegister_2_8_32_44_inst0__config_en;
  wire  ConfigRegister_2_8_32_44_inst0__reset;
  ConfigRegister_2_8_32_44 ConfigRegister_2_8_32_44_inst0(
    .O(ConfigRegister_2_8_32_44_inst0__O),
    .clk(ConfigRegister_2_8_32_44_inst0__clk),
    .config_addr(ConfigRegister_2_8_32_44_inst0__config_addr),
    .config_data(ConfigRegister_2_8_32_44_inst0__config_data),
    .config_en(ConfigRegister_2_8_32_44_inst0__config_en),
    .reset(ConfigRegister_2_8_32_44_inst0__reset)
  );

  wire [1:0] ConfigRegister_2_8_32_46_inst0__O;
  wire  ConfigRegister_2_8_32_46_inst0__clk;
  wire [7:0] ConfigRegister_2_8_32_46_inst0__config_addr;
  wire [31:0] ConfigRegister_2_8_32_46_inst0__config_data;
  wire  ConfigRegister_2_8_32_46_inst0__config_en;
  wire  ConfigRegister_2_8_32_46_inst0__reset;
  ConfigRegister_2_8_32_46 ConfigRegister_2_8_32_46_inst0(
    .O(ConfigRegister_2_8_32_46_inst0__O),
    .clk(ConfigRegister_2_8_32_46_inst0__clk),
    .config_addr(ConfigRegister_2_8_32_46_inst0__config_addr),
    .config_data(ConfigRegister_2_8_32_46_inst0__config_data),
    .config_en(ConfigRegister_2_8_32_46_inst0__config_en),
    .reset(ConfigRegister_2_8_32_46_inst0__reset)
  );

  wire [1:0] ConfigRegister_2_8_32_48_inst0__O;
  wire  ConfigRegister_2_8_32_48_inst0__clk;
  wire [7:0] ConfigRegister_2_8_32_48_inst0__config_addr;
  wire [31:0] ConfigRegister_2_8_32_48_inst0__config_data;
  wire  ConfigRegister_2_8_32_48_inst0__config_en;
  wire  ConfigRegister_2_8_32_48_inst0__reset;
  ConfigRegister_2_8_32_48 ConfigRegister_2_8_32_48_inst0(
    .O(ConfigRegister_2_8_32_48_inst0__O),
    .clk(ConfigRegister_2_8_32_48_inst0__clk),
    .config_addr(ConfigRegister_2_8_32_48_inst0__config_addr),
    .config_data(ConfigRegister_2_8_32_48_inst0__config_data),
    .config_en(ConfigRegister_2_8_32_48_inst0__config_en),
    .reset(ConfigRegister_2_8_32_48_inst0__reset)
  );

  wire [1:0] ConfigRegister_2_8_32_4_inst0__O;
  wire  ConfigRegister_2_8_32_4_inst0__clk;
  wire [7:0] ConfigRegister_2_8_32_4_inst0__config_addr;
  wire [31:0] ConfigRegister_2_8_32_4_inst0__config_data;
  wire  ConfigRegister_2_8_32_4_inst0__config_en;
  wire  ConfigRegister_2_8_32_4_inst0__reset;
  ConfigRegister_2_8_32_4 ConfigRegister_2_8_32_4_inst0(
    .O(ConfigRegister_2_8_32_4_inst0__O),
    .clk(ConfigRegister_2_8_32_4_inst0__clk),
    .config_addr(ConfigRegister_2_8_32_4_inst0__config_addr),
    .config_data(ConfigRegister_2_8_32_4_inst0__config_data),
    .config_en(ConfigRegister_2_8_32_4_inst0__config_en),
    .reset(ConfigRegister_2_8_32_4_inst0__reset)
  );

  wire [1:0] ConfigRegister_2_8_32_50_inst0__O;
  wire  ConfigRegister_2_8_32_50_inst0__clk;
  wire [7:0] ConfigRegister_2_8_32_50_inst0__config_addr;
  wire [31:0] ConfigRegister_2_8_32_50_inst0__config_data;
  wire  ConfigRegister_2_8_32_50_inst0__config_en;
  wire  ConfigRegister_2_8_32_50_inst0__reset;
  ConfigRegister_2_8_32_50 ConfigRegister_2_8_32_50_inst0(
    .O(ConfigRegister_2_8_32_50_inst0__O),
    .clk(ConfigRegister_2_8_32_50_inst0__clk),
    .config_addr(ConfigRegister_2_8_32_50_inst0__config_addr),
    .config_data(ConfigRegister_2_8_32_50_inst0__config_data),
    .config_en(ConfigRegister_2_8_32_50_inst0__config_en),
    .reset(ConfigRegister_2_8_32_50_inst0__reset)
  );

  wire [1:0] ConfigRegister_2_8_32_52_inst0__O;
  wire  ConfigRegister_2_8_32_52_inst0__clk;
  wire [7:0] ConfigRegister_2_8_32_52_inst0__config_addr;
  wire [31:0] ConfigRegister_2_8_32_52_inst0__config_data;
  wire  ConfigRegister_2_8_32_52_inst0__config_en;
  wire  ConfigRegister_2_8_32_52_inst0__reset;
  ConfigRegister_2_8_32_52 ConfigRegister_2_8_32_52_inst0(
    .O(ConfigRegister_2_8_32_52_inst0__O),
    .clk(ConfigRegister_2_8_32_52_inst0__clk),
    .config_addr(ConfigRegister_2_8_32_52_inst0__config_addr),
    .config_data(ConfigRegister_2_8_32_52_inst0__config_data),
    .config_en(ConfigRegister_2_8_32_52_inst0__config_en),
    .reset(ConfigRegister_2_8_32_52_inst0__reset)
  );

  wire [1:0] ConfigRegister_2_8_32_54_inst0__O;
  wire  ConfigRegister_2_8_32_54_inst0__clk;
  wire [7:0] ConfigRegister_2_8_32_54_inst0__config_addr;
  wire [31:0] ConfigRegister_2_8_32_54_inst0__config_data;
  wire  ConfigRegister_2_8_32_54_inst0__config_en;
  wire  ConfigRegister_2_8_32_54_inst0__reset;
  ConfigRegister_2_8_32_54 ConfigRegister_2_8_32_54_inst0(
    .O(ConfigRegister_2_8_32_54_inst0__O),
    .clk(ConfigRegister_2_8_32_54_inst0__clk),
    .config_addr(ConfigRegister_2_8_32_54_inst0__config_addr),
    .config_data(ConfigRegister_2_8_32_54_inst0__config_data),
    .config_en(ConfigRegister_2_8_32_54_inst0__config_en),
    .reset(ConfigRegister_2_8_32_54_inst0__reset)
  );

  wire [1:0] ConfigRegister_2_8_32_56_inst0__O;
  wire  ConfigRegister_2_8_32_56_inst0__clk;
  wire [7:0] ConfigRegister_2_8_32_56_inst0__config_addr;
  wire [31:0] ConfigRegister_2_8_32_56_inst0__config_data;
  wire  ConfigRegister_2_8_32_56_inst0__config_en;
  wire  ConfigRegister_2_8_32_56_inst0__reset;
  ConfigRegister_2_8_32_56 ConfigRegister_2_8_32_56_inst0(
    .O(ConfigRegister_2_8_32_56_inst0__O),
    .clk(ConfigRegister_2_8_32_56_inst0__clk),
    .config_addr(ConfigRegister_2_8_32_56_inst0__config_addr),
    .config_data(ConfigRegister_2_8_32_56_inst0__config_data),
    .config_en(ConfigRegister_2_8_32_56_inst0__config_en),
    .reset(ConfigRegister_2_8_32_56_inst0__reset)
  );

  wire [1:0] ConfigRegister_2_8_32_58_inst0__O;
  wire  ConfigRegister_2_8_32_58_inst0__clk;
  wire [7:0] ConfigRegister_2_8_32_58_inst0__config_addr;
  wire [31:0] ConfigRegister_2_8_32_58_inst0__config_data;
  wire  ConfigRegister_2_8_32_58_inst0__config_en;
  wire  ConfigRegister_2_8_32_58_inst0__reset;
  ConfigRegister_2_8_32_58 ConfigRegister_2_8_32_58_inst0(
    .O(ConfigRegister_2_8_32_58_inst0__O),
    .clk(ConfigRegister_2_8_32_58_inst0__clk),
    .config_addr(ConfigRegister_2_8_32_58_inst0__config_addr),
    .config_data(ConfigRegister_2_8_32_58_inst0__config_data),
    .config_en(ConfigRegister_2_8_32_58_inst0__config_en),
    .reset(ConfigRegister_2_8_32_58_inst0__reset)
  );

  wire [1:0] ConfigRegister_2_8_32_60_inst0__O;
  wire  ConfigRegister_2_8_32_60_inst0__clk;
  wire [7:0] ConfigRegister_2_8_32_60_inst0__config_addr;
  wire [31:0] ConfigRegister_2_8_32_60_inst0__config_data;
  wire  ConfigRegister_2_8_32_60_inst0__config_en;
  wire  ConfigRegister_2_8_32_60_inst0__reset;
  ConfigRegister_2_8_32_60 ConfigRegister_2_8_32_60_inst0(
    .O(ConfigRegister_2_8_32_60_inst0__O),
    .clk(ConfigRegister_2_8_32_60_inst0__clk),
    .config_addr(ConfigRegister_2_8_32_60_inst0__config_addr),
    .config_data(ConfigRegister_2_8_32_60_inst0__config_data),
    .config_en(ConfigRegister_2_8_32_60_inst0__config_en),
    .reset(ConfigRegister_2_8_32_60_inst0__reset)
  );

  wire [1:0] ConfigRegister_2_8_32_62_inst0__O;
  wire  ConfigRegister_2_8_32_62_inst0__clk;
  wire [7:0] ConfigRegister_2_8_32_62_inst0__config_addr;
  wire [31:0] ConfigRegister_2_8_32_62_inst0__config_data;
  wire  ConfigRegister_2_8_32_62_inst0__config_en;
  wire  ConfigRegister_2_8_32_62_inst0__reset;
  ConfigRegister_2_8_32_62 ConfigRegister_2_8_32_62_inst0(
    .O(ConfigRegister_2_8_32_62_inst0__O),
    .clk(ConfigRegister_2_8_32_62_inst0__clk),
    .config_addr(ConfigRegister_2_8_32_62_inst0__config_addr),
    .config_data(ConfigRegister_2_8_32_62_inst0__config_data),
    .config_en(ConfigRegister_2_8_32_62_inst0__config_en),
    .reset(ConfigRegister_2_8_32_62_inst0__reset)
  );

  wire [1:0] ConfigRegister_2_8_32_64_inst0__O;
  wire  ConfigRegister_2_8_32_64_inst0__clk;
  wire [7:0] ConfigRegister_2_8_32_64_inst0__config_addr;
  wire [31:0] ConfigRegister_2_8_32_64_inst0__config_data;
  wire  ConfigRegister_2_8_32_64_inst0__config_en;
  wire  ConfigRegister_2_8_32_64_inst0__reset;
  ConfigRegister_2_8_32_64 ConfigRegister_2_8_32_64_inst0(
    .O(ConfigRegister_2_8_32_64_inst0__O),
    .clk(ConfigRegister_2_8_32_64_inst0__clk),
    .config_addr(ConfigRegister_2_8_32_64_inst0__config_addr),
    .config_data(ConfigRegister_2_8_32_64_inst0__config_data),
    .config_en(ConfigRegister_2_8_32_64_inst0__config_en),
    .reset(ConfigRegister_2_8_32_64_inst0__reset)
  );

  wire [1:0] ConfigRegister_2_8_32_66_inst0__O;
  wire  ConfigRegister_2_8_32_66_inst0__clk;
  wire [7:0] ConfigRegister_2_8_32_66_inst0__config_addr;
  wire [31:0] ConfigRegister_2_8_32_66_inst0__config_data;
  wire  ConfigRegister_2_8_32_66_inst0__config_en;
  wire  ConfigRegister_2_8_32_66_inst0__reset;
  ConfigRegister_2_8_32_66 ConfigRegister_2_8_32_66_inst0(
    .O(ConfigRegister_2_8_32_66_inst0__O),
    .clk(ConfigRegister_2_8_32_66_inst0__clk),
    .config_addr(ConfigRegister_2_8_32_66_inst0__config_addr),
    .config_data(ConfigRegister_2_8_32_66_inst0__config_data),
    .config_en(ConfigRegister_2_8_32_66_inst0__config_en),
    .reset(ConfigRegister_2_8_32_66_inst0__reset)
  );

  wire [1:0] ConfigRegister_2_8_32_68_inst0__O;
  wire  ConfigRegister_2_8_32_68_inst0__clk;
  wire [7:0] ConfigRegister_2_8_32_68_inst0__config_addr;
  wire [31:0] ConfigRegister_2_8_32_68_inst0__config_data;
  wire  ConfigRegister_2_8_32_68_inst0__config_en;
  wire  ConfigRegister_2_8_32_68_inst0__reset;
  ConfigRegister_2_8_32_68 ConfigRegister_2_8_32_68_inst0(
    .O(ConfigRegister_2_8_32_68_inst0__O),
    .clk(ConfigRegister_2_8_32_68_inst0__clk),
    .config_addr(ConfigRegister_2_8_32_68_inst0__config_addr),
    .config_data(ConfigRegister_2_8_32_68_inst0__config_data),
    .config_en(ConfigRegister_2_8_32_68_inst0__config_en),
    .reset(ConfigRegister_2_8_32_68_inst0__reset)
  );

  wire [1:0] ConfigRegister_2_8_32_6_inst0__O;
  wire  ConfigRegister_2_8_32_6_inst0__clk;
  wire [7:0] ConfigRegister_2_8_32_6_inst0__config_addr;
  wire [31:0] ConfigRegister_2_8_32_6_inst0__config_data;
  wire  ConfigRegister_2_8_32_6_inst0__config_en;
  wire  ConfigRegister_2_8_32_6_inst0__reset;
  ConfigRegister_2_8_32_6 ConfigRegister_2_8_32_6_inst0(
    .O(ConfigRegister_2_8_32_6_inst0__O),
    .clk(ConfigRegister_2_8_32_6_inst0__clk),
    .config_addr(ConfigRegister_2_8_32_6_inst0__config_addr),
    .config_data(ConfigRegister_2_8_32_6_inst0__config_data),
    .config_en(ConfigRegister_2_8_32_6_inst0__config_en),
    .reset(ConfigRegister_2_8_32_6_inst0__reset)
  );

  wire [1:0] ConfigRegister_2_8_32_70_inst0__O;
  wire  ConfigRegister_2_8_32_70_inst0__clk;
  wire [7:0] ConfigRegister_2_8_32_70_inst0__config_addr;
  wire [31:0] ConfigRegister_2_8_32_70_inst0__config_data;
  wire  ConfigRegister_2_8_32_70_inst0__config_en;
  wire  ConfigRegister_2_8_32_70_inst0__reset;
  ConfigRegister_2_8_32_70 ConfigRegister_2_8_32_70_inst0(
    .O(ConfigRegister_2_8_32_70_inst0__O),
    .clk(ConfigRegister_2_8_32_70_inst0__clk),
    .config_addr(ConfigRegister_2_8_32_70_inst0__config_addr),
    .config_data(ConfigRegister_2_8_32_70_inst0__config_data),
    .config_en(ConfigRegister_2_8_32_70_inst0__config_en),
    .reset(ConfigRegister_2_8_32_70_inst0__reset)
  );

  wire [1:0] ConfigRegister_2_8_32_72_inst0__O;
  wire  ConfigRegister_2_8_32_72_inst0__clk;
  wire [7:0] ConfigRegister_2_8_32_72_inst0__config_addr;
  wire [31:0] ConfigRegister_2_8_32_72_inst0__config_data;
  wire  ConfigRegister_2_8_32_72_inst0__config_en;
  wire  ConfigRegister_2_8_32_72_inst0__reset;
  ConfigRegister_2_8_32_72 ConfigRegister_2_8_32_72_inst0(
    .O(ConfigRegister_2_8_32_72_inst0__O),
    .clk(ConfigRegister_2_8_32_72_inst0__clk),
    .config_addr(ConfigRegister_2_8_32_72_inst0__config_addr),
    .config_data(ConfigRegister_2_8_32_72_inst0__config_data),
    .config_en(ConfigRegister_2_8_32_72_inst0__config_en),
    .reset(ConfigRegister_2_8_32_72_inst0__reset)
  );

  wire [1:0] ConfigRegister_2_8_32_74_inst0__O;
  wire  ConfigRegister_2_8_32_74_inst0__clk;
  wire [7:0] ConfigRegister_2_8_32_74_inst0__config_addr;
  wire [31:0] ConfigRegister_2_8_32_74_inst0__config_data;
  wire  ConfigRegister_2_8_32_74_inst0__config_en;
  wire  ConfigRegister_2_8_32_74_inst0__reset;
  ConfigRegister_2_8_32_74 ConfigRegister_2_8_32_74_inst0(
    .O(ConfigRegister_2_8_32_74_inst0__O),
    .clk(ConfigRegister_2_8_32_74_inst0__clk),
    .config_addr(ConfigRegister_2_8_32_74_inst0__config_addr),
    .config_data(ConfigRegister_2_8_32_74_inst0__config_data),
    .config_en(ConfigRegister_2_8_32_74_inst0__config_en),
    .reset(ConfigRegister_2_8_32_74_inst0__reset)
  );

  wire [1:0] ConfigRegister_2_8_32_76_inst0__O;
  wire  ConfigRegister_2_8_32_76_inst0__clk;
  wire [7:0] ConfigRegister_2_8_32_76_inst0__config_addr;
  wire [31:0] ConfigRegister_2_8_32_76_inst0__config_data;
  wire  ConfigRegister_2_8_32_76_inst0__config_en;
  wire  ConfigRegister_2_8_32_76_inst0__reset;
  ConfigRegister_2_8_32_76 ConfigRegister_2_8_32_76_inst0(
    .O(ConfigRegister_2_8_32_76_inst0__O),
    .clk(ConfigRegister_2_8_32_76_inst0__clk),
    .config_addr(ConfigRegister_2_8_32_76_inst0__config_addr),
    .config_data(ConfigRegister_2_8_32_76_inst0__config_data),
    .config_en(ConfigRegister_2_8_32_76_inst0__config_en),
    .reset(ConfigRegister_2_8_32_76_inst0__reset)
  );

  wire [1:0] ConfigRegister_2_8_32_78_inst0__O;
  wire  ConfigRegister_2_8_32_78_inst0__clk;
  wire [7:0] ConfigRegister_2_8_32_78_inst0__config_addr;
  wire [31:0] ConfigRegister_2_8_32_78_inst0__config_data;
  wire  ConfigRegister_2_8_32_78_inst0__config_en;
  wire  ConfigRegister_2_8_32_78_inst0__reset;
  ConfigRegister_2_8_32_78 ConfigRegister_2_8_32_78_inst0(
    .O(ConfigRegister_2_8_32_78_inst0__O),
    .clk(ConfigRegister_2_8_32_78_inst0__clk),
    .config_addr(ConfigRegister_2_8_32_78_inst0__config_addr),
    .config_data(ConfigRegister_2_8_32_78_inst0__config_data),
    .config_en(ConfigRegister_2_8_32_78_inst0__config_en),
    .reset(ConfigRegister_2_8_32_78_inst0__reset)
  );

  wire [1:0] ConfigRegister_2_8_32_8_inst0__O;
  wire  ConfigRegister_2_8_32_8_inst0__clk;
  wire [7:0] ConfigRegister_2_8_32_8_inst0__config_addr;
  wire [31:0] ConfigRegister_2_8_32_8_inst0__config_data;
  wire  ConfigRegister_2_8_32_8_inst0__config_en;
  wire  ConfigRegister_2_8_32_8_inst0__reset;
  ConfigRegister_2_8_32_8 ConfigRegister_2_8_32_8_inst0(
    .O(ConfigRegister_2_8_32_8_inst0__O),
    .clk(ConfigRegister_2_8_32_8_inst0__clk),
    .config_addr(ConfigRegister_2_8_32_8_inst0__config_addr),
    .config_data(ConfigRegister_2_8_32_8_inst0__config_data),
    .config_en(ConfigRegister_2_8_32_8_inst0__config_en),
    .reset(ConfigRegister_2_8_32_8_inst0__reset)
  );

  wire [15:0] MuxWrapper_2_16_inst0__I_0;
  wire [15:0] MuxWrapper_2_16_inst0__I_1;
  wire [15:0] MuxWrapper_2_16_inst0__O;
  wire [0:0] MuxWrapper_2_16_inst0__S;
  MuxWrapper_2_16 MuxWrapper_2_16_inst0(
    .I_0(MuxWrapper_2_16_inst0__I_0),
    .I_1(MuxWrapper_2_16_inst0__I_1),
    .O(MuxWrapper_2_16_inst0__O),
    .S(MuxWrapper_2_16_inst0__S)
  );

  wire [15:0] MuxWrapper_2_16_inst1__I_0;
  wire [15:0] MuxWrapper_2_16_inst1__I_1;
  wire [15:0] MuxWrapper_2_16_inst1__O;
  wire [0:0] MuxWrapper_2_16_inst1__S;
  MuxWrapper_2_16 MuxWrapper_2_16_inst1(
    .I_0(MuxWrapper_2_16_inst1__I_0),
    .I_1(MuxWrapper_2_16_inst1__I_1),
    .O(MuxWrapper_2_16_inst1__O),
    .S(MuxWrapper_2_16_inst1__S)
  );

  wire [15:0] MuxWrapper_2_16_inst10__I_0;
  wire [15:0] MuxWrapper_2_16_inst10__I_1;
  wire [15:0] MuxWrapper_2_16_inst10__O;
  wire [0:0] MuxWrapper_2_16_inst10__S;
  MuxWrapper_2_16 MuxWrapper_2_16_inst10(
    .I_0(MuxWrapper_2_16_inst10__I_0),
    .I_1(MuxWrapper_2_16_inst10__I_1),
    .O(MuxWrapper_2_16_inst10__O),
    .S(MuxWrapper_2_16_inst10__S)
  );

  wire [15:0] MuxWrapper_2_16_inst11__I_0;
  wire [15:0] MuxWrapper_2_16_inst11__I_1;
  wire [15:0] MuxWrapper_2_16_inst11__O;
  wire [0:0] MuxWrapper_2_16_inst11__S;
  MuxWrapper_2_16 MuxWrapper_2_16_inst11(
    .I_0(MuxWrapper_2_16_inst11__I_0),
    .I_1(MuxWrapper_2_16_inst11__I_1),
    .O(MuxWrapper_2_16_inst11__O),
    .S(MuxWrapper_2_16_inst11__S)
  );

  wire [15:0] MuxWrapper_2_16_inst12__I_0;
  wire [15:0] MuxWrapper_2_16_inst12__I_1;
  wire [15:0] MuxWrapper_2_16_inst12__O;
  wire [0:0] MuxWrapper_2_16_inst12__S;
  MuxWrapper_2_16 MuxWrapper_2_16_inst12(
    .I_0(MuxWrapper_2_16_inst12__I_0),
    .I_1(MuxWrapper_2_16_inst12__I_1),
    .O(MuxWrapper_2_16_inst12__O),
    .S(MuxWrapper_2_16_inst12__S)
  );

  wire [15:0] MuxWrapper_2_16_inst13__I_0;
  wire [15:0] MuxWrapper_2_16_inst13__I_1;
  wire [15:0] MuxWrapper_2_16_inst13__O;
  wire [0:0] MuxWrapper_2_16_inst13__S;
  MuxWrapper_2_16 MuxWrapper_2_16_inst13(
    .I_0(MuxWrapper_2_16_inst13__I_0),
    .I_1(MuxWrapper_2_16_inst13__I_1),
    .O(MuxWrapper_2_16_inst13__O),
    .S(MuxWrapper_2_16_inst13__S)
  );

  wire [15:0] MuxWrapper_2_16_inst14__I_0;
  wire [15:0] MuxWrapper_2_16_inst14__I_1;
  wire [15:0] MuxWrapper_2_16_inst14__O;
  wire [0:0] MuxWrapper_2_16_inst14__S;
  MuxWrapper_2_16 MuxWrapper_2_16_inst14(
    .I_0(MuxWrapper_2_16_inst14__I_0),
    .I_1(MuxWrapper_2_16_inst14__I_1),
    .O(MuxWrapper_2_16_inst14__O),
    .S(MuxWrapper_2_16_inst14__S)
  );

  wire [15:0] MuxWrapper_2_16_inst15__I_0;
  wire [15:0] MuxWrapper_2_16_inst15__I_1;
  wire [15:0] MuxWrapper_2_16_inst15__O;
  wire [0:0] MuxWrapper_2_16_inst15__S;
  MuxWrapper_2_16 MuxWrapper_2_16_inst15(
    .I_0(MuxWrapper_2_16_inst15__I_0),
    .I_1(MuxWrapper_2_16_inst15__I_1),
    .O(MuxWrapper_2_16_inst15__O),
    .S(MuxWrapper_2_16_inst15__S)
  );

  wire [15:0] MuxWrapper_2_16_inst16__I_0;
  wire [15:0] MuxWrapper_2_16_inst16__I_1;
  wire [15:0] MuxWrapper_2_16_inst16__O;
  wire [0:0] MuxWrapper_2_16_inst16__S;
  MuxWrapper_2_16 MuxWrapper_2_16_inst16(
    .I_0(MuxWrapper_2_16_inst16__I_0),
    .I_1(MuxWrapper_2_16_inst16__I_1),
    .O(MuxWrapper_2_16_inst16__O),
    .S(MuxWrapper_2_16_inst16__S)
  );

  wire [15:0] MuxWrapper_2_16_inst17__I_0;
  wire [15:0] MuxWrapper_2_16_inst17__I_1;
  wire [15:0] MuxWrapper_2_16_inst17__O;
  wire [0:0] MuxWrapper_2_16_inst17__S;
  MuxWrapper_2_16 MuxWrapper_2_16_inst17(
    .I_0(MuxWrapper_2_16_inst17__I_0),
    .I_1(MuxWrapper_2_16_inst17__I_1),
    .O(MuxWrapper_2_16_inst17__O),
    .S(MuxWrapper_2_16_inst17__S)
  );

  wire [15:0] MuxWrapper_2_16_inst18__I_0;
  wire [15:0] MuxWrapper_2_16_inst18__I_1;
  wire [15:0] MuxWrapper_2_16_inst18__O;
  wire [0:0] MuxWrapper_2_16_inst18__S;
  MuxWrapper_2_16 MuxWrapper_2_16_inst18(
    .I_0(MuxWrapper_2_16_inst18__I_0),
    .I_1(MuxWrapper_2_16_inst18__I_1),
    .O(MuxWrapper_2_16_inst18__O),
    .S(MuxWrapper_2_16_inst18__S)
  );

  wire [15:0] MuxWrapper_2_16_inst19__I_0;
  wire [15:0] MuxWrapper_2_16_inst19__I_1;
  wire [15:0] MuxWrapper_2_16_inst19__O;
  wire [0:0] MuxWrapper_2_16_inst19__S;
  MuxWrapper_2_16 MuxWrapper_2_16_inst19(
    .I_0(MuxWrapper_2_16_inst19__I_0),
    .I_1(MuxWrapper_2_16_inst19__I_1),
    .O(MuxWrapper_2_16_inst19__O),
    .S(MuxWrapper_2_16_inst19__S)
  );

  wire [15:0] MuxWrapper_2_16_inst2__I_0;
  wire [15:0] MuxWrapper_2_16_inst2__I_1;
  wire [15:0] MuxWrapper_2_16_inst2__O;
  wire [0:0] MuxWrapper_2_16_inst2__S;
  MuxWrapper_2_16 MuxWrapper_2_16_inst2(
    .I_0(MuxWrapper_2_16_inst2__I_0),
    .I_1(MuxWrapper_2_16_inst2__I_1),
    .O(MuxWrapper_2_16_inst2__O),
    .S(MuxWrapper_2_16_inst2__S)
  );

  wire [15:0] MuxWrapper_2_16_inst3__I_0;
  wire [15:0] MuxWrapper_2_16_inst3__I_1;
  wire [15:0] MuxWrapper_2_16_inst3__O;
  wire [0:0] MuxWrapper_2_16_inst3__S;
  MuxWrapper_2_16 MuxWrapper_2_16_inst3(
    .I_0(MuxWrapper_2_16_inst3__I_0),
    .I_1(MuxWrapper_2_16_inst3__I_1),
    .O(MuxWrapper_2_16_inst3__O),
    .S(MuxWrapper_2_16_inst3__S)
  );

  wire [15:0] MuxWrapper_2_16_inst4__I_0;
  wire [15:0] MuxWrapper_2_16_inst4__I_1;
  wire [15:0] MuxWrapper_2_16_inst4__O;
  wire [0:0] MuxWrapper_2_16_inst4__S;
  MuxWrapper_2_16 MuxWrapper_2_16_inst4(
    .I_0(MuxWrapper_2_16_inst4__I_0),
    .I_1(MuxWrapper_2_16_inst4__I_1),
    .O(MuxWrapper_2_16_inst4__O),
    .S(MuxWrapper_2_16_inst4__S)
  );

  wire [15:0] MuxWrapper_2_16_inst5__I_0;
  wire [15:0] MuxWrapper_2_16_inst5__I_1;
  wire [15:0] MuxWrapper_2_16_inst5__O;
  wire [0:0] MuxWrapper_2_16_inst5__S;
  MuxWrapper_2_16 MuxWrapper_2_16_inst5(
    .I_0(MuxWrapper_2_16_inst5__I_0),
    .I_1(MuxWrapper_2_16_inst5__I_1),
    .O(MuxWrapper_2_16_inst5__O),
    .S(MuxWrapper_2_16_inst5__S)
  );

  wire [15:0] MuxWrapper_2_16_inst6__I_0;
  wire [15:0] MuxWrapper_2_16_inst6__I_1;
  wire [15:0] MuxWrapper_2_16_inst6__O;
  wire [0:0] MuxWrapper_2_16_inst6__S;
  MuxWrapper_2_16 MuxWrapper_2_16_inst6(
    .I_0(MuxWrapper_2_16_inst6__I_0),
    .I_1(MuxWrapper_2_16_inst6__I_1),
    .O(MuxWrapper_2_16_inst6__O),
    .S(MuxWrapper_2_16_inst6__S)
  );

  wire [15:0] MuxWrapper_2_16_inst7__I_0;
  wire [15:0] MuxWrapper_2_16_inst7__I_1;
  wire [15:0] MuxWrapper_2_16_inst7__O;
  wire [0:0] MuxWrapper_2_16_inst7__S;
  MuxWrapper_2_16 MuxWrapper_2_16_inst7(
    .I_0(MuxWrapper_2_16_inst7__I_0),
    .I_1(MuxWrapper_2_16_inst7__I_1),
    .O(MuxWrapper_2_16_inst7__O),
    .S(MuxWrapper_2_16_inst7__S)
  );

  wire [15:0] MuxWrapper_2_16_inst8__I_0;
  wire [15:0] MuxWrapper_2_16_inst8__I_1;
  wire [15:0] MuxWrapper_2_16_inst8__O;
  wire [0:0] MuxWrapper_2_16_inst8__S;
  MuxWrapper_2_16 MuxWrapper_2_16_inst8(
    .I_0(MuxWrapper_2_16_inst8__I_0),
    .I_1(MuxWrapper_2_16_inst8__I_1),
    .O(MuxWrapper_2_16_inst8__O),
    .S(MuxWrapper_2_16_inst8__S)
  );

  wire [15:0] MuxWrapper_2_16_inst9__I_0;
  wire [15:0] MuxWrapper_2_16_inst9__I_1;
  wire [15:0] MuxWrapper_2_16_inst9__O;
  wire [0:0] MuxWrapper_2_16_inst9__S;
  MuxWrapper_2_16 MuxWrapper_2_16_inst9(
    .I_0(MuxWrapper_2_16_inst9__I_0),
    .I_1(MuxWrapper_2_16_inst9__I_1),
    .O(MuxWrapper_2_16_inst9__O),
    .S(MuxWrapper_2_16_inst9__S)
  );

  wire [0:0] MuxWrapper_2_1_inst0__I_0;
  wire [0:0] MuxWrapper_2_1_inst0__I_1;
  wire [0:0] MuxWrapper_2_1_inst0__O;
  wire [0:0] MuxWrapper_2_1_inst0__S;
  MuxWrapper_2_1 MuxWrapper_2_1_inst0(
    .I_0(MuxWrapper_2_1_inst0__I_0),
    .I_1(MuxWrapper_2_1_inst0__I_1),
    .O(MuxWrapper_2_1_inst0__O),
    .S(MuxWrapper_2_1_inst0__S)
  );

  wire [0:0] MuxWrapper_2_1_inst1__I_0;
  wire [0:0] MuxWrapper_2_1_inst1__I_1;
  wire [0:0] MuxWrapper_2_1_inst1__O;
  wire [0:0] MuxWrapper_2_1_inst1__S;
  MuxWrapper_2_1 MuxWrapper_2_1_inst1(
    .I_0(MuxWrapper_2_1_inst1__I_0),
    .I_1(MuxWrapper_2_1_inst1__I_1),
    .O(MuxWrapper_2_1_inst1__O),
    .S(MuxWrapper_2_1_inst1__S)
  );

  wire [0:0] MuxWrapper_2_1_inst10__I_0;
  wire [0:0] MuxWrapper_2_1_inst10__I_1;
  wire [0:0] MuxWrapper_2_1_inst10__O;
  wire [0:0] MuxWrapper_2_1_inst10__S;
  MuxWrapper_2_1 MuxWrapper_2_1_inst10(
    .I_0(MuxWrapper_2_1_inst10__I_0),
    .I_1(MuxWrapper_2_1_inst10__I_1),
    .O(MuxWrapper_2_1_inst10__O),
    .S(MuxWrapper_2_1_inst10__S)
  );

  wire [0:0] MuxWrapper_2_1_inst11__I_0;
  wire [0:0] MuxWrapper_2_1_inst11__I_1;
  wire [0:0] MuxWrapper_2_1_inst11__O;
  wire [0:0] MuxWrapper_2_1_inst11__S;
  MuxWrapper_2_1 MuxWrapper_2_1_inst11(
    .I_0(MuxWrapper_2_1_inst11__I_0),
    .I_1(MuxWrapper_2_1_inst11__I_1),
    .O(MuxWrapper_2_1_inst11__O),
    .S(MuxWrapper_2_1_inst11__S)
  );

  wire [0:0] MuxWrapper_2_1_inst12__I_0;
  wire [0:0] MuxWrapper_2_1_inst12__I_1;
  wire [0:0] MuxWrapper_2_1_inst12__O;
  wire [0:0] MuxWrapper_2_1_inst12__S;
  MuxWrapper_2_1 MuxWrapper_2_1_inst12(
    .I_0(MuxWrapper_2_1_inst12__I_0),
    .I_1(MuxWrapper_2_1_inst12__I_1),
    .O(MuxWrapper_2_1_inst12__O),
    .S(MuxWrapper_2_1_inst12__S)
  );

  wire [0:0] MuxWrapper_2_1_inst13__I_0;
  wire [0:0] MuxWrapper_2_1_inst13__I_1;
  wire [0:0] MuxWrapper_2_1_inst13__O;
  wire [0:0] MuxWrapper_2_1_inst13__S;
  MuxWrapper_2_1 MuxWrapper_2_1_inst13(
    .I_0(MuxWrapper_2_1_inst13__I_0),
    .I_1(MuxWrapper_2_1_inst13__I_1),
    .O(MuxWrapper_2_1_inst13__O),
    .S(MuxWrapper_2_1_inst13__S)
  );

  wire [0:0] MuxWrapper_2_1_inst14__I_0;
  wire [0:0] MuxWrapper_2_1_inst14__I_1;
  wire [0:0] MuxWrapper_2_1_inst14__O;
  wire [0:0] MuxWrapper_2_1_inst14__S;
  MuxWrapper_2_1 MuxWrapper_2_1_inst14(
    .I_0(MuxWrapper_2_1_inst14__I_0),
    .I_1(MuxWrapper_2_1_inst14__I_1),
    .O(MuxWrapper_2_1_inst14__O),
    .S(MuxWrapper_2_1_inst14__S)
  );

  wire [0:0] MuxWrapper_2_1_inst15__I_0;
  wire [0:0] MuxWrapper_2_1_inst15__I_1;
  wire [0:0] MuxWrapper_2_1_inst15__O;
  wire [0:0] MuxWrapper_2_1_inst15__S;
  MuxWrapper_2_1 MuxWrapper_2_1_inst15(
    .I_0(MuxWrapper_2_1_inst15__I_0),
    .I_1(MuxWrapper_2_1_inst15__I_1),
    .O(MuxWrapper_2_1_inst15__O),
    .S(MuxWrapper_2_1_inst15__S)
  );

  wire [0:0] MuxWrapper_2_1_inst16__I_0;
  wire [0:0] MuxWrapper_2_1_inst16__I_1;
  wire [0:0] MuxWrapper_2_1_inst16__O;
  wire [0:0] MuxWrapper_2_1_inst16__S;
  MuxWrapper_2_1 MuxWrapper_2_1_inst16(
    .I_0(MuxWrapper_2_1_inst16__I_0),
    .I_1(MuxWrapper_2_1_inst16__I_1),
    .O(MuxWrapper_2_1_inst16__O),
    .S(MuxWrapper_2_1_inst16__S)
  );

  wire [0:0] MuxWrapper_2_1_inst17__I_0;
  wire [0:0] MuxWrapper_2_1_inst17__I_1;
  wire [0:0] MuxWrapper_2_1_inst17__O;
  wire [0:0] MuxWrapper_2_1_inst17__S;
  MuxWrapper_2_1 MuxWrapper_2_1_inst17(
    .I_0(MuxWrapper_2_1_inst17__I_0),
    .I_1(MuxWrapper_2_1_inst17__I_1),
    .O(MuxWrapper_2_1_inst17__O),
    .S(MuxWrapper_2_1_inst17__S)
  );

  wire [0:0] MuxWrapper_2_1_inst18__I_0;
  wire [0:0] MuxWrapper_2_1_inst18__I_1;
  wire [0:0] MuxWrapper_2_1_inst18__O;
  wire [0:0] MuxWrapper_2_1_inst18__S;
  MuxWrapper_2_1 MuxWrapper_2_1_inst18(
    .I_0(MuxWrapper_2_1_inst18__I_0),
    .I_1(MuxWrapper_2_1_inst18__I_1),
    .O(MuxWrapper_2_1_inst18__O),
    .S(MuxWrapper_2_1_inst18__S)
  );

  wire [0:0] MuxWrapper_2_1_inst19__I_0;
  wire [0:0] MuxWrapper_2_1_inst19__I_1;
  wire [0:0] MuxWrapper_2_1_inst19__O;
  wire [0:0] MuxWrapper_2_1_inst19__S;
  MuxWrapper_2_1 MuxWrapper_2_1_inst19(
    .I_0(MuxWrapper_2_1_inst19__I_0),
    .I_1(MuxWrapper_2_1_inst19__I_1),
    .O(MuxWrapper_2_1_inst19__O),
    .S(MuxWrapper_2_1_inst19__S)
  );

  wire [0:0] MuxWrapper_2_1_inst2__I_0;
  wire [0:0] MuxWrapper_2_1_inst2__I_1;
  wire [0:0] MuxWrapper_2_1_inst2__O;
  wire [0:0] MuxWrapper_2_1_inst2__S;
  MuxWrapper_2_1 MuxWrapper_2_1_inst2(
    .I_0(MuxWrapper_2_1_inst2__I_0),
    .I_1(MuxWrapper_2_1_inst2__I_1),
    .O(MuxWrapper_2_1_inst2__O),
    .S(MuxWrapper_2_1_inst2__S)
  );

  wire [0:0] MuxWrapper_2_1_inst3__I_0;
  wire [0:0] MuxWrapper_2_1_inst3__I_1;
  wire [0:0] MuxWrapper_2_1_inst3__O;
  wire [0:0] MuxWrapper_2_1_inst3__S;
  MuxWrapper_2_1 MuxWrapper_2_1_inst3(
    .I_0(MuxWrapper_2_1_inst3__I_0),
    .I_1(MuxWrapper_2_1_inst3__I_1),
    .O(MuxWrapper_2_1_inst3__O),
    .S(MuxWrapper_2_1_inst3__S)
  );

  wire [0:0] MuxWrapper_2_1_inst4__I_0;
  wire [0:0] MuxWrapper_2_1_inst4__I_1;
  wire [0:0] MuxWrapper_2_1_inst4__O;
  wire [0:0] MuxWrapper_2_1_inst4__S;
  MuxWrapper_2_1 MuxWrapper_2_1_inst4(
    .I_0(MuxWrapper_2_1_inst4__I_0),
    .I_1(MuxWrapper_2_1_inst4__I_1),
    .O(MuxWrapper_2_1_inst4__O),
    .S(MuxWrapper_2_1_inst4__S)
  );

  wire [0:0] MuxWrapper_2_1_inst5__I_0;
  wire [0:0] MuxWrapper_2_1_inst5__I_1;
  wire [0:0] MuxWrapper_2_1_inst5__O;
  wire [0:0] MuxWrapper_2_1_inst5__S;
  MuxWrapper_2_1 MuxWrapper_2_1_inst5(
    .I_0(MuxWrapper_2_1_inst5__I_0),
    .I_1(MuxWrapper_2_1_inst5__I_1),
    .O(MuxWrapper_2_1_inst5__O),
    .S(MuxWrapper_2_1_inst5__S)
  );

  wire [0:0] MuxWrapper_2_1_inst6__I_0;
  wire [0:0] MuxWrapper_2_1_inst6__I_1;
  wire [0:0] MuxWrapper_2_1_inst6__O;
  wire [0:0] MuxWrapper_2_1_inst6__S;
  MuxWrapper_2_1 MuxWrapper_2_1_inst6(
    .I_0(MuxWrapper_2_1_inst6__I_0),
    .I_1(MuxWrapper_2_1_inst6__I_1),
    .O(MuxWrapper_2_1_inst6__O),
    .S(MuxWrapper_2_1_inst6__S)
  );

  wire [0:0] MuxWrapper_2_1_inst7__I_0;
  wire [0:0] MuxWrapper_2_1_inst7__I_1;
  wire [0:0] MuxWrapper_2_1_inst7__O;
  wire [0:0] MuxWrapper_2_1_inst7__S;
  MuxWrapper_2_1 MuxWrapper_2_1_inst7(
    .I_0(MuxWrapper_2_1_inst7__I_0),
    .I_1(MuxWrapper_2_1_inst7__I_1),
    .O(MuxWrapper_2_1_inst7__O),
    .S(MuxWrapper_2_1_inst7__S)
  );

  wire [0:0] MuxWrapper_2_1_inst8__I_0;
  wire [0:0] MuxWrapper_2_1_inst8__I_1;
  wire [0:0] MuxWrapper_2_1_inst8__O;
  wire [0:0] MuxWrapper_2_1_inst8__S;
  MuxWrapper_2_1 MuxWrapper_2_1_inst8(
    .I_0(MuxWrapper_2_1_inst8__I_0),
    .I_1(MuxWrapper_2_1_inst8__I_1),
    .O(MuxWrapper_2_1_inst8__O),
    .S(MuxWrapper_2_1_inst8__S)
  );

  wire [0:0] MuxWrapper_2_1_inst9__I_0;
  wire [0:0] MuxWrapper_2_1_inst9__I_1;
  wire [0:0] MuxWrapper_2_1_inst9__O;
  wire [0:0] MuxWrapper_2_1_inst9__S;
  MuxWrapper_2_1 MuxWrapper_2_1_inst9(
    .I_0(MuxWrapper_2_1_inst9__I_0),
    .I_1(MuxWrapper_2_1_inst9__I_1),
    .O(MuxWrapper_2_1_inst9__O),
    .S(MuxWrapper_2_1_inst9__S)
  );

  wire [15:0] MuxWrapper_4_16_inst0__I_0;
  wire [15:0] MuxWrapper_4_16_inst0__I_1;
  wire [15:0] MuxWrapper_4_16_inst0__I_2;
  wire [15:0] MuxWrapper_4_16_inst0__I_3;
  wire [15:0] MuxWrapper_4_16_inst0__O;
  wire [1:0] MuxWrapper_4_16_inst0__S;
  MuxWrapper_4_16 MuxWrapper_4_16_inst0(
    .I_0(MuxWrapper_4_16_inst0__I_0),
    .I_1(MuxWrapper_4_16_inst0__I_1),
    .I_2(MuxWrapper_4_16_inst0__I_2),
    .I_3(MuxWrapper_4_16_inst0__I_3),
    .O(MuxWrapper_4_16_inst0__O),
    .S(MuxWrapper_4_16_inst0__S)
  );

  wire [15:0] MuxWrapper_4_16_inst1__I_0;
  wire [15:0] MuxWrapper_4_16_inst1__I_1;
  wire [15:0] MuxWrapper_4_16_inst1__I_2;
  wire [15:0] MuxWrapper_4_16_inst1__I_3;
  wire [15:0] MuxWrapper_4_16_inst1__O;
  wire [1:0] MuxWrapper_4_16_inst1__S;
  MuxWrapper_4_16 MuxWrapper_4_16_inst1(
    .I_0(MuxWrapper_4_16_inst1__I_0),
    .I_1(MuxWrapper_4_16_inst1__I_1),
    .I_2(MuxWrapper_4_16_inst1__I_2),
    .I_3(MuxWrapper_4_16_inst1__I_3),
    .O(MuxWrapper_4_16_inst1__O),
    .S(MuxWrapper_4_16_inst1__S)
  );

  wire [15:0] MuxWrapper_4_16_inst10__I_0;
  wire [15:0] MuxWrapper_4_16_inst10__I_1;
  wire [15:0] MuxWrapper_4_16_inst10__I_2;
  wire [15:0] MuxWrapper_4_16_inst10__I_3;
  wire [15:0] MuxWrapper_4_16_inst10__O;
  wire [1:0] MuxWrapper_4_16_inst10__S;
  MuxWrapper_4_16 MuxWrapper_4_16_inst10(
    .I_0(MuxWrapper_4_16_inst10__I_0),
    .I_1(MuxWrapper_4_16_inst10__I_1),
    .I_2(MuxWrapper_4_16_inst10__I_2),
    .I_3(MuxWrapper_4_16_inst10__I_3),
    .O(MuxWrapper_4_16_inst10__O),
    .S(MuxWrapper_4_16_inst10__S)
  );

  wire [15:0] MuxWrapper_4_16_inst11__I_0;
  wire [15:0] MuxWrapper_4_16_inst11__I_1;
  wire [15:0] MuxWrapper_4_16_inst11__I_2;
  wire [15:0] MuxWrapper_4_16_inst11__I_3;
  wire [15:0] MuxWrapper_4_16_inst11__O;
  wire [1:0] MuxWrapper_4_16_inst11__S;
  MuxWrapper_4_16 MuxWrapper_4_16_inst11(
    .I_0(MuxWrapper_4_16_inst11__I_0),
    .I_1(MuxWrapper_4_16_inst11__I_1),
    .I_2(MuxWrapper_4_16_inst11__I_2),
    .I_3(MuxWrapper_4_16_inst11__I_3),
    .O(MuxWrapper_4_16_inst11__O),
    .S(MuxWrapper_4_16_inst11__S)
  );

  wire [15:0] MuxWrapper_4_16_inst12__I_0;
  wire [15:0] MuxWrapper_4_16_inst12__I_1;
  wire [15:0] MuxWrapper_4_16_inst12__I_2;
  wire [15:0] MuxWrapper_4_16_inst12__I_3;
  wire [15:0] MuxWrapper_4_16_inst12__O;
  wire [1:0] MuxWrapper_4_16_inst12__S;
  MuxWrapper_4_16 MuxWrapper_4_16_inst12(
    .I_0(MuxWrapper_4_16_inst12__I_0),
    .I_1(MuxWrapper_4_16_inst12__I_1),
    .I_2(MuxWrapper_4_16_inst12__I_2),
    .I_3(MuxWrapper_4_16_inst12__I_3),
    .O(MuxWrapper_4_16_inst12__O),
    .S(MuxWrapper_4_16_inst12__S)
  );

  wire [15:0] MuxWrapper_4_16_inst13__I_0;
  wire [15:0] MuxWrapper_4_16_inst13__I_1;
  wire [15:0] MuxWrapper_4_16_inst13__I_2;
  wire [15:0] MuxWrapper_4_16_inst13__I_3;
  wire [15:0] MuxWrapper_4_16_inst13__O;
  wire [1:0] MuxWrapper_4_16_inst13__S;
  MuxWrapper_4_16 MuxWrapper_4_16_inst13(
    .I_0(MuxWrapper_4_16_inst13__I_0),
    .I_1(MuxWrapper_4_16_inst13__I_1),
    .I_2(MuxWrapper_4_16_inst13__I_2),
    .I_3(MuxWrapper_4_16_inst13__I_3),
    .O(MuxWrapper_4_16_inst13__O),
    .S(MuxWrapper_4_16_inst13__S)
  );

  wire [15:0] MuxWrapper_4_16_inst14__I_0;
  wire [15:0] MuxWrapper_4_16_inst14__I_1;
  wire [15:0] MuxWrapper_4_16_inst14__I_2;
  wire [15:0] MuxWrapper_4_16_inst14__I_3;
  wire [15:0] MuxWrapper_4_16_inst14__O;
  wire [1:0] MuxWrapper_4_16_inst14__S;
  MuxWrapper_4_16 MuxWrapper_4_16_inst14(
    .I_0(MuxWrapper_4_16_inst14__I_0),
    .I_1(MuxWrapper_4_16_inst14__I_1),
    .I_2(MuxWrapper_4_16_inst14__I_2),
    .I_3(MuxWrapper_4_16_inst14__I_3),
    .O(MuxWrapper_4_16_inst14__O),
    .S(MuxWrapper_4_16_inst14__S)
  );

  wire [15:0] MuxWrapper_4_16_inst15__I_0;
  wire [15:0] MuxWrapper_4_16_inst15__I_1;
  wire [15:0] MuxWrapper_4_16_inst15__I_2;
  wire [15:0] MuxWrapper_4_16_inst15__I_3;
  wire [15:0] MuxWrapper_4_16_inst15__O;
  wire [1:0] MuxWrapper_4_16_inst15__S;
  MuxWrapper_4_16 MuxWrapper_4_16_inst15(
    .I_0(MuxWrapper_4_16_inst15__I_0),
    .I_1(MuxWrapper_4_16_inst15__I_1),
    .I_2(MuxWrapper_4_16_inst15__I_2),
    .I_3(MuxWrapper_4_16_inst15__I_3),
    .O(MuxWrapper_4_16_inst15__O),
    .S(MuxWrapper_4_16_inst15__S)
  );

  wire [15:0] MuxWrapper_4_16_inst16__I_0;
  wire [15:0] MuxWrapper_4_16_inst16__I_1;
  wire [15:0] MuxWrapper_4_16_inst16__I_2;
  wire [15:0] MuxWrapper_4_16_inst16__I_3;
  wire [15:0] MuxWrapper_4_16_inst16__O;
  wire [1:0] MuxWrapper_4_16_inst16__S;
  MuxWrapper_4_16 MuxWrapper_4_16_inst16(
    .I_0(MuxWrapper_4_16_inst16__I_0),
    .I_1(MuxWrapper_4_16_inst16__I_1),
    .I_2(MuxWrapper_4_16_inst16__I_2),
    .I_3(MuxWrapper_4_16_inst16__I_3),
    .O(MuxWrapper_4_16_inst16__O),
    .S(MuxWrapper_4_16_inst16__S)
  );

  wire [15:0] MuxWrapper_4_16_inst17__I_0;
  wire [15:0] MuxWrapper_4_16_inst17__I_1;
  wire [15:0] MuxWrapper_4_16_inst17__I_2;
  wire [15:0] MuxWrapper_4_16_inst17__I_3;
  wire [15:0] MuxWrapper_4_16_inst17__O;
  wire [1:0] MuxWrapper_4_16_inst17__S;
  MuxWrapper_4_16 MuxWrapper_4_16_inst17(
    .I_0(MuxWrapper_4_16_inst17__I_0),
    .I_1(MuxWrapper_4_16_inst17__I_1),
    .I_2(MuxWrapper_4_16_inst17__I_2),
    .I_3(MuxWrapper_4_16_inst17__I_3),
    .O(MuxWrapper_4_16_inst17__O),
    .S(MuxWrapper_4_16_inst17__S)
  );

  wire [15:0] MuxWrapper_4_16_inst18__I_0;
  wire [15:0] MuxWrapper_4_16_inst18__I_1;
  wire [15:0] MuxWrapper_4_16_inst18__I_2;
  wire [15:0] MuxWrapper_4_16_inst18__I_3;
  wire [15:0] MuxWrapper_4_16_inst18__O;
  wire [1:0] MuxWrapper_4_16_inst18__S;
  MuxWrapper_4_16 MuxWrapper_4_16_inst18(
    .I_0(MuxWrapper_4_16_inst18__I_0),
    .I_1(MuxWrapper_4_16_inst18__I_1),
    .I_2(MuxWrapper_4_16_inst18__I_2),
    .I_3(MuxWrapper_4_16_inst18__I_3),
    .O(MuxWrapper_4_16_inst18__O),
    .S(MuxWrapper_4_16_inst18__S)
  );

  wire [15:0] MuxWrapper_4_16_inst19__I_0;
  wire [15:0] MuxWrapper_4_16_inst19__I_1;
  wire [15:0] MuxWrapper_4_16_inst19__I_2;
  wire [15:0] MuxWrapper_4_16_inst19__I_3;
  wire [15:0] MuxWrapper_4_16_inst19__O;
  wire [1:0] MuxWrapper_4_16_inst19__S;
  MuxWrapper_4_16 MuxWrapper_4_16_inst19(
    .I_0(MuxWrapper_4_16_inst19__I_0),
    .I_1(MuxWrapper_4_16_inst19__I_1),
    .I_2(MuxWrapper_4_16_inst19__I_2),
    .I_3(MuxWrapper_4_16_inst19__I_3),
    .O(MuxWrapper_4_16_inst19__O),
    .S(MuxWrapper_4_16_inst19__S)
  );

  wire [15:0] MuxWrapper_4_16_inst2__I_0;
  wire [15:0] MuxWrapper_4_16_inst2__I_1;
  wire [15:0] MuxWrapper_4_16_inst2__I_2;
  wire [15:0] MuxWrapper_4_16_inst2__I_3;
  wire [15:0] MuxWrapper_4_16_inst2__O;
  wire [1:0] MuxWrapper_4_16_inst2__S;
  MuxWrapper_4_16 MuxWrapper_4_16_inst2(
    .I_0(MuxWrapper_4_16_inst2__I_0),
    .I_1(MuxWrapper_4_16_inst2__I_1),
    .I_2(MuxWrapper_4_16_inst2__I_2),
    .I_3(MuxWrapper_4_16_inst2__I_3),
    .O(MuxWrapper_4_16_inst2__O),
    .S(MuxWrapper_4_16_inst2__S)
  );

  wire [15:0] MuxWrapper_4_16_inst3__I_0;
  wire [15:0] MuxWrapper_4_16_inst3__I_1;
  wire [15:0] MuxWrapper_4_16_inst3__I_2;
  wire [15:0] MuxWrapper_4_16_inst3__I_3;
  wire [15:0] MuxWrapper_4_16_inst3__O;
  wire [1:0] MuxWrapper_4_16_inst3__S;
  MuxWrapper_4_16 MuxWrapper_4_16_inst3(
    .I_0(MuxWrapper_4_16_inst3__I_0),
    .I_1(MuxWrapper_4_16_inst3__I_1),
    .I_2(MuxWrapper_4_16_inst3__I_2),
    .I_3(MuxWrapper_4_16_inst3__I_3),
    .O(MuxWrapper_4_16_inst3__O),
    .S(MuxWrapper_4_16_inst3__S)
  );

  wire [15:0] MuxWrapper_4_16_inst4__I_0;
  wire [15:0] MuxWrapper_4_16_inst4__I_1;
  wire [15:0] MuxWrapper_4_16_inst4__I_2;
  wire [15:0] MuxWrapper_4_16_inst4__I_3;
  wire [15:0] MuxWrapper_4_16_inst4__O;
  wire [1:0] MuxWrapper_4_16_inst4__S;
  MuxWrapper_4_16 MuxWrapper_4_16_inst4(
    .I_0(MuxWrapper_4_16_inst4__I_0),
    .I_1(MuxWrapper_4_16_inst4__I_1),
    .I_2(MuxWrapper_4_16_inst4__I_2),
    .I_3(MuxWrapper_4_16_inst4__I_3),
    .O(MuxWrapper_4_16_inst4__O),
    .S(MuxWrapper_4_16_inst4__S)
  );

  wire [15:0] MuxWrapper_4_16_inst5__I_0;
  wire [15:0] MuxWrapper_4_16_inst5__I_1;
  wire [15:0] MuxWrapper_4_16_inst5__I_2;
  wire [15:0] MuxWrapper_4_16_inst5__I_3;
  wire [15:0] MuxWrapper_4_16_inst5__O;
  wire [1:0] MuxWrapper_4_16_inst5__S;
  MuxWrapper_4_16 MuxWrapper_4_16_inst5(
    .I_0(MuxWrapper_4_16_inst5__I_0),
    .I_1(MuxWrapper_4_16_inst5__I_1),
    .I_2(MuxWrapper_4_16_inst5__I_2),
    .I_3(MuxWrapper_4_16_inst5__I_3),
    .O(MuxWrapper_4_16_inst5__O),
    .S(MuxWrapper_4_16_inst5__S)
  );

  wire [15:0] MuxWrapper_4_16_inst6__I_0;
  wire [15:0] MuxWrapper_4_16_inst6__I_1;
  wire [15:0] MuxWrapper_4_16_inst6__I_2;
  wire [15:0] MuxWrapper_4_16_inst6__I_3;
  wire [15:0] MuxWrapper_4_16_inst6__O;
  wire [1:0] MuxWrapper_4_16_inst6__S;
  MuxWrapper_4_16 MuxWrapper_4_16_inst6(
    .I_0(MuxWrapper_4_16_inst6__I_0),
    .I_1(MuxWrapper_4_16_inst6__I_1),
    .I_2(MuxWrapper_4_16_inst6__I_2),
    .I_3(MuxWrapper_4_16_inst6__I_3),
    .O(MuxWrapper_4_16_inst6__O),
    .S(MuxWrapper_4_16_inst6__S)
  );

  wire [15:0] MuxWrapper_4_16_inst7__I_0;
  wire [15:0] MuxWrapper_4_16_inst7__I_1;
  wire [15:0] MuxWrapper_4_16_inst7__I_2;
  wire [15:0] MuxWrapper_4_16_inst7__I_3;
  wire [15:0] MuxWrapper_4_16_inst7__O;
  wire [1:0] MuxWrapper_4_16_inst7__S;
  MuxWrapper_4_16 MuxWrapper_4_16_inst7(
    .I_0(MuxWrapper_4_16_inst7__I_0),
    .I_1(MuxWrapper_4_16_inst7__I_1),
    .I_2(MuxWrapper_4_16_inst7__I_2),
    .I_3(MuxWrapper_4_16_inst7__I_3),
    .O(MuxWrapper_4_16_inst7__O),
    .S(MuxWrapper_4_16_inst7__S)
  );

  wire [15:0] MuxWrapper_4_16_inst8__I_0;
  wire [15:0] MuxWrapper_4_16_inst8__I_1;
  wire [15:0] MuxWrapper_4_16_inst8__I_2;
  wire [15:0] MuxWrapper_4_16_inst8__I_3;
  wire [15:0] MuxWrapper_4_16_inst8__O;
  wire [1:0] MuxWrapper_4_16_inst8__S;
  MuxWrapper_4_16 MuxWrapper_4_16_inst8(
    .I_0(MuxWrapper_4_16_inst8__I_0),
    .I_1(MuxWrapper_4_16_inst8__I_1),
    .I_2(MuxWrapper_4_16_inst8__I_2),
    .I_3(MuxWrapper_4_16_inst8__I_3),
    .O(MuxWrapper_4_16_inst8__O),
    .S(MuxWrapper_4_16_inst8__S)
  );

  wire [15:0] MuxWrapper_4_16_inst9__I_0;
  wire [15:0] MuxWrapper_4_16_inst9__I_1;
  wire [15:0] MuxWrapper_4_16_inst9__I_2;
  wire [15:0] MuxWrapper_4_16_inst9__I_3;
  wire [15:0] MuxWrapper_4_16_inst9__O;
  wire [1:0] MuxWrapper_4_16_inst9__S;
  MuxWrapper_4_16 MuxWrapper_4_16_inst9(
    .I_0(MuxWrapper_4_16_inst9__I_0),
    .I_1(MuxWrapper_4_16_inst9__I_1),
    .I_2(MuxWrapper_4_16_inst9__I_2),
    .I_3(MuxWrapper_4_16_inst9__I_3),
    .O(MuxWrapper_4_16_inst9__O),
    .S(MuxWrapper_4_16_inst9__S)
  );

  wire [0:0] MuxWrapper_4_1_inst0__I_0;
  wire [0:0] MuxWrapper_4_1_inst0__I_1;
  wire [0:0] MuxWrapper_4_1_inst0__I_2;
  wire [0:0] MuxWrapper_4_1_inst0__I_3;
  wire [0:0] MuxWrapper_4_1_inst0__O;
  wire [1:0] MuxWrapper_4_1_inst0__S;
  MuxWrapper_4_1 MuxWrapper_4_1_inst0(
    .I_0(MuxWrapper_4_1_inst0__I_0),
    .I_1(MuxWrapper_4_1_inst0__I_1),
    .I_2(MuxWrapper_4_1_inst0__I_2),
    .I_3(MuxWrapper_4_1_inst0__I_3),
    .O(MuxWrapper_4_1_inst0__O),
    .S(MuxWrapper_4_1_inst0__S)
  );

  wire [0:0] MuxWrapper_4_1_inst1__I_0;
  wire [0:0] MuxWrapper_4_1_inst1__I_1;
  wire [0:0] MuxWrapper_4_1_inst1__I_2;
  wire [0:0] MuxWrapper_4_1_inst1__I_3;
  wire [0:0] MuxWrapper_4_1_inst1__O;
  wire [1:0] MuxWrapper_4_1_inst1__S;
  MuxWrapper_4_1 MuxWrapper_4_1_inst1(
    .I_0(MuxWrapper_4_1_inst1__I_0),
    .I_1(MuxWrapper_4_1_inst1__I_1),
    .I_2(MuxWrapper_4_1_inst1__I_2),
    .I_3(MuxWrapper_4_1_inst1__I_3),
    .O(MuxWrapper_4_1_inst1__O),
    .S(MuxWrapper_4_1_inst1__S)
  );

  wire [0:0] MuxWrapper_4_1_inst10__I_0;
  wire [0:0] MuxWrapper_4_1_inst10__I_1;
  wire [0:0] MuxWrapper_4_1_inst10__I_2;
  wire [0:0] MuxWrapper_4_1_inst10__I_3;
  wire [0:0] MuxWrapper_4_1_inst10__O;
  wire [1:0] MuxWrapper_4_1_inst10__S;
  MuxWrapper_4_1 MuxWrapper_4_1_inst10(
    .I_0(MuxWrapper_4_1_inst10__I_0),
    .I_1(MuxWrapper_4_1_inst10__I_1),
    .I_2(MuxWrapper_4_1_inst10__I_2),
    .I_3(MuxWrapper_4_1_inst10__I_3),
    .O(MuxWrapper_4_1_inst10__O),
    .S(MuxWrapper_4_1_inst10__S)
  );

  wire [0:0] MuxWrapper_4_1_inst11__I_0;
  wire [0:0] MuxWrapper_4_1_inst11__I_1;
  wire [0:0] MuxWrapper_4_1_inst11__I_2;
  wire [0:0] MuxWrapper_4_1_inst11__I_3;
  wire [0:0] MuxWrapper_4_1_inst11__O;
  wire [1:0] MuxWrapper_4_1_inst11__S;
  MuxWrapper_4_1 MuxWrapper_4_1_inst11(
    .I_0(MuxWrapper_4_1_inst11__I_0),
    .I_1(MuxWrapper_4_1_inst11__I_1),
    .I_2(MuxWrapper_4_1_inst11__I_2),
    .I_3(MuxWrapper_4_1_inst11__I_3),
    .O(MuxWrapper_4_1_inst11__O),
    .S(MuxWrapper_4_1_inst11__S)
  );

  wire [0:0] MuxWrapper_4_1_inst12__I_0;
  wire [0:0] MuxWrapper_4_1_inst12__I_1;
  wire [0:0] MuxWrapper_4_1_inst12__I_2;
  wire [0:0] MuxWrapper_4_1_inst12__I_3;
  wire [0:0] MuxWrapper_4_1_inst12__O;
  wire [1:0] MuxWrapper_4_1_inst12__S;
  MuxWrapper_4_1 MuxWrapper_4_1_inst12(
    .I_0(MuxWrapper_4_1_inst12__I_0),
    .I_1(MuxWrapper_4_1_inst12__I_1),
    .I_2(MuxWrapper_4_1_inst12__I_2),
    .I_3(MuxWrapper_4_1_inst12__I_3),
    .O(MuxWrapper_4_1_inst12__O),
    .S(MuxWrapper_4_1_inst12__S)
  );

  wire [0:0] MuxWrapper_4_1_inst13__I_0;
  wire [0:0] MuxWrapper_4_1_inst13__I_1;
  wire [0:0] MuxWrapper_4_1_inst13__I_2;
  wire [0:0] MuxWrapper_4_1_inst13__I_3;
  wire [0:0] MuxWrapper_4_1_inst13__O;
  wire [1:0] MuxWrapper_4_1_inst13__S;
  MuxWrapper_4_1 MuxWrapper_4_1_inst13(
    .I_0(MuxWrapper_4_1_inst13__I_0),
    .I_1(MuxWrapper_4_1_inst13__I_1),
    .I_2(MuxWrapper_4_1_inst13__I_2),
    .I_3(MuxWrapper_4_1_inst13__I_3),
    .O(MuxWrapper_4_1_inst13__O),
    .S(MuxWrapper_4_1_inst13__S)
  );

  wire [0:0] MuxWrapper_4_1_inst14__I_0;
  wire [0:0] MuxWrapper_4_1_inst14__I_1;
  wire [0:0] MuxWrapper_4_1_inst14__I_2;
  wire [0:0] MuxWrapper_4_1_inst14__I_3;
  wire [0:0] MuxWrapper_4_1_inst14__O;
  wire [1:0] MuxWrapper_4_1_inst14__S;
  MuxWrapper_4_1 MuxWrapper_4_1_inst14(
    .I_0(MuxWrapper_4_1_inst14__I_0),
    .I_1(MuxWrapper_4_1_inst14__I_1),
    .I_2(MuxWrapper_4_1_inst14__I_2),
    .I_3(MuxWrapper_4_1_inst14__I_3),
    .O(MuxWrapper_4_1_inst14__O),
    .S(MuxWrapper_4_1_inst14__S)
  );

  wire [0:0] MuxWrapper_4_1_inst15__I_0;
  wire [0:0] MuxWrapper_4_1_inst15__I_1;
  wire [0:0] MuxWrapper_4_1_inst15__I_2;
  wire [0:0] MuxWrapper_4_1_inst15__I_3;
  wire [0:0] MuxWrapper_4_1_inst15__O;
  wire [1:0] MuxWrapper_4_1_inst15__S;
  MuxWrapper_4_1 MuxWrapper_4_1_inst15(
    .I_0(MuxWrapper_4_1_inst15__I_0),
    .I_1(MuxWrapper_4_1_inst15__I_1),
    .I_2(MuxWrapper_4_1_inst15__I_2),
    .I_3(MuxWrapper_4_1_inst15__I_3),
    .O(MuxWrapper_4_1_inst15__O),
    .S(MuxWrapper_4_1_inst15__S)
  );

  wire [0:0] MuxWrapper_4_1_inst16__I_0;
  wire [0:0] MuxWrapper_4_1_inst16__I_1;
  wire [0:0] MuxWrapper_4_1_inst16__I_2;
  wire [0:0] MuxWrapper_4_1_inst16__I_3;
  wire [0:0] MuxWrapper_4_1_inst16__O;
  wire [1:0] MuxWrapper_4_1_inst16__S;
  MuxWrapper_4_1 MuxWrapper_4_1_inst16(
    .I_0(MuxWrapper_4_1_inst16__I_0),
    .I_1(MuxWrapper_4_1_inst16__I_1),
    .I_2(MuxWrapper_4_1_inst16__I_2),
    .I_3(MuxWrapper_4_1_inst16__I_3),
    .O(MuxWrapper_4_1_inst16__O),
    .S(MuxWrapper_4_1_inst16__S)
  );

  wire [0:0] MuxWrapper_4_1_inst17__I_0;
  wire [0:0] MuxWrapper_4_1_inst17__I_1;
  wire [0:0] MuxWrapper_4_1_inst17__I_2;
  wire [0:0] MuxWrapper_4_1_inst17__I_3;
  wire [0:0] MuxWrapper_4_1_inst17__O;
  wire [1:0] MuxWrapper_4_1_inst17__S;
  MuxWrapper_4_1 MuxWrapper_4_1_inst17(
    .I_0(MuxWrapper_4_1_inst17__I_0),
    .I_1(MuxWrapper_4_1_inst17__I_1),
    .I_2(MuxWrapper_4_1_inst17__I_2),
    .I_3(MuxWrapper_4_1_inst17__I_3),
    .O(MuxWrapper_4_1_inst17__O),
    .S(MuxWrapper_4_1_inst17__S)
  );

  wire [0:0] MuxWrapper_4_1_inst18__I_0;
  wire [0:0] MuxWrapper_4_1_inst18__I_1;
  wire [0:0] MuxWrapper_4_1_inst18__I_2;
  wire [0:0] MuxWrapper_4_1_inst18__I_3;
  wire [0:0] MuxWrapper_4_1_inst18__O;
  wire [1:0] MuxWrapper_4_1_inst18__S;
  MuxWrapper_4_1 MuxWrapper_4_1_inst18(
    .I_0(MuxWrapper_4_1_inst18__I_0),
    .I_1(MuxWrapper_4_1_inst18__I_1),
    .I_2(MuxWrapper_4_1_inst18__I_2),
    .I_3(MuxWrapper_4_1_inst18__I_3),
    .O(MuxWrapper_4_1_inst18__O),
    .S(MuxWrapper_4_1_inst18__S)
  );

  wire [0:0] MuxWrapper_4_1_inst19__I_0;
  wire [0:0] MuxWrapper_4_1_inst19__I_1;
  wire [0:0] MuxWrapper_4_1_inst19__I_2;
  wire [0:0] MuxWrapper_4_1_inst19__I_3;
  wire [0:0] MuxWrapper_4_1_inst19__O;
  wire [1:0] MuxWrapper_4_1_inst19__S;
  MuxWrapper_4_1 MuxWrapper_4_1_inst19(
    .I_0(MuxWrapper_4_1_inst19__I_0),
    .I_1(MuxWrapper_4_1_inst19__I_1),
    .I_2(MuxWrapper_4_1_inst19__I_2),
    .I_3(MuxWrapper_4_1_inst19__I_3),
    .O(MuxWrapper_4_1_inst19__O),
    .S(MuxWrapper_4_1_inst19__S)
  );

  wire [0:0] MuxWrapper_4_1_inst2__I_0;
  wire [0:0] MuxWrapper_4_1_inst2__I_1;
  wire [0:0] MuxWrapper_4_1_inst2__I_2;
  wire [0:0] MuxWrapper_4_1_inst2__I_3;
  wire [0:0] MuxWrapper_4_1_inst2__O;
  wire [1:0] MuxWrapper_4_1_inst2__S;
  MuxWrapper_4_1 MuxWrapper_4_1_inst2(
    .I_0(MuxWrapper_4_1_inst2__I_0),
    .I_1(MuxWrapper_4_1_inst2__I_1),
    .I_2(MuxWrapper_4_1_inst2__I_2),
    .I_3(MuxWrapper_4_1_inst2__I_3),
    .O(MuxWrapper_4_1_inst2__O),
    .S(MuxWrapper_4_1_inst2__S)
  );

  wire [0:0] MuxWrapper_4_1_inst3__I_0;
  wire [0:0] MuxWrapper_4_1_inst3__I_1;
  wire [0:0] MuxWrapper_4_1_inst3__I_2;
  wire [0:0] MuxWrapper_4_1_inst3__I_3;
  wire [0:0] MuxWrapper_4_1_inst3__O;
  wire [1:0] MuxWrapper_4_1_inst3__S;
  MuxWrapper_4_1 MuxWrapper_4_1_inst3(
    .I_0(MuxWrapper_4_1_inst3__I_0),
    .I_1(MuxWrapper_4_1_inst3__I_1),
    .I_2(MuxWrapper_4_1_inst3__I_2),
    .I_3(MuxWrapper_4_1_inst3__I_3),
    .O(MuxWrapper_4_1_inst3__O),
    .S(MuxWrapper_4_1_inst3__S)
  );

  wire [0:0] MuxWrapper_4_1_inst4__I_0;
  wire [0:0] MuxWrapper_4_1_inst4__I_1;
  wire [0:0] MuxWrapper_4_1_inst4__I_2;
  wire [0:0] MuxWrapper_4_1_inst4__I_3;
  wire [0:0] MuxWrapper_4_1_inst4__O;
  wire [1:0] MuxWrapper_4_1_inst4__S;
  MuxWrapper_4_1 MuxWrapper_4_1_inst4(
    .I_0(MuxWrapper_4_1_inst4__I_0),
    .I_1(MuxWrapper_4_1_inst4__I_1),
    .I_2(MuxWrapper_4_1_inst4__I_2),
    .I_3(MuxWrapper_4_1_inst4__I_3),
    .O(MuxWrapper_4_1_inst4__O),
    .S(MuxWrapper_4_1_inst4__S)
  );

  wire [0:0] MuxWrapper_4_1_inst5__I_0;
  wire [0:0] MuxWrapper_4_1_inst5__I_1;
  wire [0:0] MuxWrapper_4_1_inst5__I_2;
  wire [0:0] MuxWrapper_4_1_inst5__I_3;
  wire [0:0] MuxWrapper_4_1_inst5__O;
  wire [1:0] MuxWrapper_4_1_inst5__S;
  MuxWrapper_4_1 MuxWrapper_4_1_inst5(
    .I_0(MuxWrapper_4_1_inst5__I_0),
    .I_1(MuxWrapper_4_1_inst5__I_1),
    .I_2(MuxWrapper_4_1_inst5__I_2),
    .I_3(MuxWrapper_4_1_inst5__I_3),
    .O(MuxWrapper_4_1_inst5__O),
    .S(MuxWrapper_4_1_inst5__S)
  );

  wire [0:0] MuxWrapper_4_1_inst6__I_0;
  wire [0:0] MuxWrapper_4_1_inst6__I_1;
  wire [0:0] MuxWrapper_4_1_inst6__I_2;
  wire [0:0] MuxWrapper_4_1_inst6__I_3;
  wire [0:0] MuxWrapper_4_1_inst6__O;
  wire [1:0] MuxWrapper_4_1_inst6__S;
  MuxWrapper_4_1 MuxWrapper_4_1_inst6(
    .I_0(MuxWrapper_4_1_inst6__I_0),
    .I_1(MuxWrapper_4_1_inst6__I_1),
    .I_2(MuxWrapper_4_1_inst6__I_2),
    .I_3(MuxWrapper_4_1_inst6__I_3),
    .O(MuxWrapper_4_1_inst6__O),
    .S(MuxWrapper_4_1_inst6__S)
  );

  wire [0:0] MuxWrapper_4_1_inst7__I_0;
  wire [0:0] MuxWrapper_4_1_inst7__I_1;
  wire [0:0] MuxWrapper_4_1_inst7__I_2;
  wire [0:0] MuxWrapper_4_1_inst7__I_3;
  wire [0:0] MuxWrapper_4_1_inst7__O;
  wire [1:0] MuxWrapper_4_1_inst7__S;
  MuxWrapper_4_1 MuxWrapper_4_1_inst7(
    .I_0(MuxWrapper_4_1_inst7__I_0),
    .I_1(MuxWrapper_4_1_inst7__I_1),
    .I_2(MuxWrapper_4_1_inst7__I_2),
    .I_3(MuxWrapper_4_1_inst7__I_3),
    .O(MuxWrapper_4_1_inst7__O),
    .S(MuxWrapper_4_1_inst7__S)
  );

  wire [0:0] MuxWrapper_4_1_inst8__I_0;
  wire [0:0] MuxWrapper_4_1_inst8__I_1;
  wire [0:0] MuxWrapper_4_1_inst8__I_2;
  wire [0:0] MuxWrapper_4_1_inst8__I_3;
  wire [0:0] MuxWrapper_4_1_inst8__O;
  wire [1:0] MuxWrapper_4_1_inst8__S;
  MuxWrapper_4_1 MuxWrapper_4_1_inst8(
    .I_0(MuxWrapper_4_1_inst8__I_0),
    .I_1(MuxWrapper_4_1_inst8__I_1),
    .I_2(MuxWrapper_4_1_inst8__I_2),
    .I_3(MuxWrapper_4_1_inst8__I_3),
    .O(MuxWrapper_4_1_inst8__O),
    .S(MuxWrapper_4_1_inst8__S)
  );

  wire [0:0] MuxWrapper_4_1_inst9__I_0;
  wire [0:0] MuxWrapper_4_1_inst9__I_1;
  wire [0:0] MuxWrapper_4_1_inst9__I_2;
  wire [0:0] MuxWrapper_4_1_inst9__I_3;
  wire [0:0] MuxWrapper_4_1_inst9__O;
  wire [1:0] MuxWrapper_4_1_inst9__S;
  MuxWrapper_4_1 MuxWrapper_4_1_inst9(
    .I_0(MuxWrapper_4_1_inst9__I_0),
    .I_1(MuxWrapper_4_1_inst9__I_1),
    .I_2(MuxWrapper_4_1_inst9__I_2),
    .I_3(MuxWrapper_4_1_inst9__I_3),
    .O(MuxWrapper_4_1_inst9__O),
    .S(MuxWrapper_4_1_inst9__S)
  );

  wire [31:0] MuxWrapper_80_32_inst0__I_0;
  wire [31:0] MuxWrapper_80_32_inst0__I_1;
  wire [31:0] MuxWrapper_80_32_inst0__I_10;
  wire [31:0] MuxWrapper_80_32_inst0__I_11;
  wire [31:0] MuxWrapper_80_32_inst0__I_12;
  wire [31:0] MuxWrapper_80_32_inst0__I_13;
  wire [31:0] MuxWrapper_80_32_inst0__I_14;
  wire [31:0] MuxWrapper_80_32_inst0__I_15;
  wire [31:0] MuxWrapper_80_32_inst0__I_16;
  wire [31:0] MuxWrapper_80_32_inst0__I_17;
  wire [31:0] MuxWrapper_80_32_inst0__I_18;
  wire [31:0] MuxWrapper_80_32_inst0__I_19;
  wire [31:0] MuxWrapper_80_32_inst0__I_2;
  wire [31:0] MuxWrapper_80_32_inst0__I_20;
  wire [31:0] MuxWrapper_80_32_inst0__I_21;
  wire [31:0] MuxWrapper_80_32_inst0__I_22;
  wire [31:0] MuxWrapper_80_32_inst0__I_23;
  wire [31:0] MuxWrapper_80_32_inst0__I_24;
  wire [31:0] MuxWrapper_80_32_inst0__I_25;
  wire [31:0] MuxWrapper_80_32_inst0__I_26;
  wire [31:0] MuxWrapper_80_32_inst0__I_27;
  wire [31:0] MuxWrapper_80_32_inst0__I_28;
  wire [31:0] MuxWrapper_80_32_inst0__I_29;
  wire [31:0] MuxWrapper_80_32_inst0__I_3;
  wire [31:0] MuxWrapper_80_32_inst0__I_30;
  wire [31:0] MuxWrapper_80_32_inst0__I_31;
  wire [31:0] MuxWrapper_80_32_inst0__I_32;
  wire [31:0] MuxWrapper_80_32_inst0__I_33;
  wire [31:0] MuxWrapper_80_32_inst0__I_34;
  wire [31:0] MuxWrapper_80_32_inst0__I_35;
  wire [31:0] MuxWrapper_80_32_inst0__I_36;
  wire [31:0] MuxWrapper_80_32_inst0__I_37;
  wire [31:0] MuxWrapper_80_32_inst0__I_38;
  wire [31:0] MuxWrapper_80_32_inst0__I_39;
  wire [31:0] MuxWrapper_80_32_inst0__I_4;
  wire [31:0] MuxWrapper_80_32_inst0__I_40;
  wire [31:0] MuxWrapper_80_32_inst0__I_41;
  wire [31:0] MuxWrapper_80_32_inst0__I_42;
  wire [31:0] MuxWrapper_80_32_inst0__I_43;
  wire [31:0] MuxWrapper_80_32_inst0__I_44;
  wire [31:0] MuxWrapper_80_32_inst0__I_45;
  wire [31:0] MuxWrapper_80_32_inst0__I_46;
  wire [31:0] MuxWrapper_80_32_inst0__I_47;
  wire [31:0] MuxWrapper_80_32_inst0__I_48;
  wire [31:0] MuxWrapper_80_32_inst0__I_49;
  wire [31:0] MuxWrapper_80_32_inst0__I_5;
  wire [31:0] MuxWrapper_80_32_inst0__I_50;
  wire [31:0] MuxWrapper_80_32_inst0__I_51;
  wire [31:0] MuxWrapper_80_32_inst0__I_52;
  wire [31:0] MuxWrapper_80_32_inst0__I_53;
  wire [31:0] MuxWrapper_80_32_inst0__I_54;
  wire [31:0] MuxWrapper_80_32_inst0__I_55;
  wire [31:0] MuxWrapper_80_32_inst0__I_56;
  wire [31:0] MuxWrapper_80_32_inst0__I_57;
  wire [31:0] MuxWrapper_80_32_inst0__I_58;
  wire [31:0] MuxWrapper_80_32_inst0__I_59;
  wire [31:0] MuxWrapper_80_32_inst0__I_6;
  wire [31:0] MuxWrapper_80_32_inst0__I_60;
  wire [31:0] MuxWrapper_80_32_inst0__I_61;
  wire [31:0] MuxWrapper_80_32_inst0__I_62;
  wire [31:0] MuxWrapper_80_32_inst0__I_63;
  wire [31:0] MuxWrapper_80_32_inst0__I_64;
  wire [31:0] MuxWrapper_80_32_inst0__I_65;
  wire [31:0] MuxWrapper_80_32_inst0__I_66;
  wire [31:0] MuxWrapper_80_32_inst0__I_67;
  wire [31:0] MuxWrapper_80_32_inst0__I_68;
  wire [31:0] MuxWrapper_80_32_inst0__I_69;
  wire [31:0] MuxWrapper_80_32_inst0__I_7;
  wire [31:0] MuxWrapper_80_32_inst0__I_70;
  wire [31:0] MuxWrapper_80_32_inst0__I_71;
  wire [31:0] MuxWrapper_80_32_inst0__I_72;
  wire [31:0] MuxWrapper_80_32_inst0__I_73;
  wire [31:0] MuxWrapper_80_32_inst0__I_74;
  wire [31:0] MuxWrapper_80_32_inst0__I_75;
  wire [31:0] MuxWrapper_80_32_inst0__I_76;
  wire [31:0] MuxWrapper_80_32_inst0__I_77;
  wire [31:0] MuxWrapper_80_32_inst0__I_78;
  wire [31:0] MuxWrapper_80_32_inst0__I_79;
  wire [31:0] MuxWrapper_80_32_inst0__I_8;
  wire [31:0] MuxWrapper_80_32_inst0__I_9;
  wire [31:0] MuxWrapper_80_32_inst0__O;
  wire [6:0] MuxWrapper_80_32_inst0__S;
  MuxWrapper_80_32 MuxWrapper_80_32_inst0(
    .I_0(MuxWrapper_80_32_inst0__I_0),
    .I_1(MuxWrapper_80_32_inst0__I_1),
    .I_10(MuxWrapper_80_32_inst0__I_10),
    .I_11(MuxWrapper_80_32_inst0__I_11),
    .I_12(MuxWrapper_80_32_inst0__I_12),
    .I_13(MuxWrapper_80_32_inst0__I_13),
    .I_14(MuxWrapper_80_32_inst0__I_14),
    .I_15(MuxWrapper_80_32_inst0__I_15),
    .I_16(MuxWrapper_80_32_inst0__I_16),
    .I_17(MuxWrapper_80_32_inst0__I_17),
    .I_18(MuxWrapper_80_32_inst0__I_18),
    .I_19(MuxWrapper_80_32_inst0__I_19),
    .I_2(MuxWrapper_80_32_inst0__I_2),
    .I_20(MuxWrapper_80_32_inst0__I_20),
    .I_21(MuxWrapper_80_32_inst0__I_21),
    .I_22(MuxWrapper_80_32_inst0__I_22),
    .I_23(MuxWrapper_80_32_inst0__I_23),
    .I_24(MuxWrapper_80_32_inst0__I_24),
    .I_25(MuxWrapper_80_32_inst0__I_25),
    .I_26(MuxWrapper_80_32_inst0__I_26),
    .I_27(MuxWrapper_80_32_inst0__I_27),
    .I_28(MuxWrapper_80_32_inst0__I_28),
    .I_29(MuxWrapper_80_32_inst0__I_29),
    .I_3(MuxWrapper_80_32_inst0__I_3),
    .I_30(MuxWrapper_80_32_inst0__I_30),
    .I_31(MuxWrapper_80_32_inst0__I_31),
    .I_32(MuxWrapper_80_32_inst0__I_32),
    .I_33(MuxWrapper_80_32_inst0__I_33),
    .I_34(MuxWrapper_80_32_inst0__I_34),
    .I_35(MuxWrapper_80_32_inst0__I_35),
    .I_36(MuxWrapper_80_32_inst0__I_36),
    .I_37(MuxWrapper_80_32_inst0__I_37),
    .I_38(MuxWrapper_80_32_inst0__I_38),
    .I_39(MuxWrapper_80_32_inst0__I_39),
    .I_4(MuxWrapper_80_32_inst0__I_4),
    .I_40(MuxWrapper_80_32_inst0__I_40),
    .I_41(MuxWrapper_80_32_inst0__I_41),
    .I_42(MuxWrapper_80_32_inst0__I_42),
    .I_43(MuxWrapper_80_32_inst0__I_43),
    .I_44(MuxWrapper_80_32_inst0__I_44),
    .I_45(MuxWrapper_80_32_inst0__I_45),
    .I_46(MuxWrapper_80_32_inst0__I_46),
    .I_47(MuxWrapper_80_32_inst0__I_47),
    .I_48(MuxWrapper_80_32_inst0__I_48),
    .I_49(MuxWrapper_80_32_inst0__I_49),
    .I_5(MuxWrapper_80_32_inst0__I_5),
    .I_50(MuxWrapper_80_32_inst0__I_50),
    .I_51(MuxWrapper_80_32_inst0__I_51),
    .I_52(MuxWrapper_80_32_inst0__I_52),
    .I_53(MuxWrapper_80_32_inst0__I_53),
    .I_54(MuxWrapper_80_32_inst0__I_54),
    .I_55(MuxWrapper_80_32_inst0__I_55),
    .I_56(MuxWrapper_80_32_inst0__I_56),
    .I_57(MuxWrapper_80_32_inst0__I_57),
    .I_58(MuxWrapper_80_32_inst0__I_58),
    .I_59(MuxWrapper_80_32_inst0__I_59),
    .I_6(MuxWrapper_80_32_inst0__I_6),
    .I_60(MuxWrapper_80_32_inst0__I_60),
    .I_61(MuxWrapper_80_32_inst0__I_61),
    .I_62(MuxWrapper_80_32_inst0__I_62),
    .I_63(MuxWrapper_80_32_inst0__I_63),
    .I_64(MuxWrapper_80_32_inst0__I_64),
    .I_65(MuxWrapper_80_32_inst0__I_65),
    .I_66(MuxWrapper_80_32_inst0__I_66),
    .I_67(MuxWrapper_80_32_inst0__I_67),
    .I_68(MuxWrapper_80_32_inst0__I_68),
    .I_69(MuxWrapper_80_32_inst0__I_69),
    .I_7(MuxWrapper_80_32_inst0__I_7),
    .I_70(MuxWrapper_80_32_inst0__I_70),
    .I_71(MuxWrapper_80_32_inst0__I_71),
    .I_72(MuxWrapper_80_32_inst0__I_72),
    .I_73(MuxWrapper_80_32_inst0__I_73),
    .I_74(MuxWrapper_80_32_inst0__I_74),
    .I_75(MuxWrapper_80_32_inst0__I_75),
    .I_76(MuxWrapper_80_32_inst0__I_76),
    .I_77(MuxWrapper_80_32_inst0__I_77),
    .I_78(MuxWrapper_80_32_inst0__I_78),
    .I_79(MuxWrapper_80_32_inst0__I_79),
    .I_8(MuxWrapper_80_32_inst0__I_8),
    .I_9(MuxWrapper_80_32_inst0__I_9),
    .O(MuxWrapper_80_32_inst0__O),
    .S(MuxWrapper_80_32_inst0__S)
  );

  wire [0:0] ZextWrapper_1_32_inst0__I;
  wire [31:0] ZextWrapper_1_32_inst0__O;
  ZextWrapper_1_32 ZextWrapper_1_32_inst0(
    .I(ZextWrapper_1_32_inst0__I),
    .O(ZextWrapper_1_32_inst0__O)
  );

  wire [0:0] ZextWrapper_1_32_inst1__I;
  wire [31:0] ZextWrapper_1_32_inst1__O;
  ZextWrapper_1_32 ZextWrapper_1_32_inst1(
    .I(ZextWrapper_1_32_inst1__I),
    .O(ZextWrapper_1_32_inst1__O)
  );

  wire [0:0] ZextWrapper_1_32_inst10__I;
  wire [31:0] ZextWrapper_1_32_inst10__O;
  ZextWrapper_1_32 ZextWrapper_1_32_inst10(
    .I(ZextWrapper_1_32_inst10__I),
    .O(ZextWrapper_1_32_inst10__O)
  );

  wire [0:0] ZextWrapper_1_32_inst11__I;
  wire [31:0] ZextWrapper_1_32_inst11__O;
  ZextWrapper_1_32 ZextWrapper_1_32_inst11(
    .I(ZextWrapper_1_32_inst11__I),
    .O(ZextWrapper_1_32_inst11__O)
  );

  wire [0:0] ZextWrapper_1_32_inst12__I;
  wire [31:0] ZextWrapper_1_32_inst12__O;
  ZextWrapper_1_32 ZextWrapper_1_32_inst12(
    .I(ZextWrapper_1_32_inst12__I),
    .O(ZextWrapper_1_32_inst12__O)
  );

  wire [0:0] ZextWrapper_1_32_inst13__I;
  wire [31:0] ZextWrapper_1_32_inst13__O;
  ZextWrapper_1_32 ZextWrapper_1_32_inst13(
    .I(ZextWrapper_1_32_inst13__I),
    .O(ZextWrapper_1_32_inst13__O)
  );

  wire [0:0] ZextWrapper_1_32_inst14__I;
  wire [31:0] ZextWrapper_1_32_inst14__O;
  ZextWrapper_1_32 ZextWrapper_1_32_inst14(
    .I(ZextWrapper_1_32_inst14__I),
    .O(ZextWrapper_1_32_inst14__O)
  );

  wire [0:0] ZextWrapper_1_32_inst15__I;
  wire [31:0] ZextWrapper_1_32_inst15__O;
  ZextWrapper_1_32 ZextWrapper_1_32_inst15(
    .I(ZextWrapper_1_32_inst15__I),
    .O(ZextWrapper_1_32_inst15__O)
  );

  wire [0:0] ZextWrapper_1_32_inst16__I;
  wire [31:0] ZextWrapper_1_32_inst16__O;
  ZextWrapper_1_32 ZextWrapper_1_32_inst16(
    .I(ZextWrapper_1_32_inst16__I),
    .O(ZextWrapper_1_32_inst16__O)
  );

  wire [0:0] ZextWrapper_1_32_inst17__I;
  wire [31:0] ZextWrapper_1_32_inst17__O;
  ZextWrapper_1_32 ZextWrapper_1_32_inst17(
    .I(ZextWrapper_1_32_inst17__I),
    .O(ZextWrapper_1_32_inst17__O)
  );

  wire [0:0] ZextWrapper_1_32_inst18__I;
  wire [31:0] ZextWrapper_1_32_inst18__O;
  ZextWrapper_1_32 ZextWrapper_1_32_inst18(
    .I(ZextWrapper_1_32_inst18__I),
    .O(ZextWrapper_1_32_inst18__O)
  );

  wire [0:0] ZextWrapper_1_32_inst19__I;
  wire [31:0] ZextWrapper_1_32_inst19__O;
  ZextWrapper_1_32 ZextWrapper_1_32_inst19(
    .I(ZextWrapper_1_32_inst19__I),
    .O(ZextWrapper_1_32_inst19__O)
  );

  wire [0:0] ZextWrapper_1_32_inst2__I;
  wire [31:0] ZextWrapper_1_32_inst2__O;
  ZextWrapper_1_32 ZextWrapper_1_32_inst2(
    .I(ZextWrapper_1_32_inst2__I),
    .O(ZextWrapper_1_32_inst2__O)
  );

  wire [0:0] ZextWrapper_1_32_inst20__I;
  wire [31:0] ZextWrapper_1_32_inst20__O;
  ZextWrapper_1_32 ZextWrapper_1_32_inst20(
    .I(ZextWrapper_1_32_inst20__I),
    .O(ZextWrapper_1_32_inst20__O)
  );

  wire [0:0] ZextWrapper_1_32_inst21__I;
  wire [31:0] ZextWrapper_1_32_inst21__O;
  ZextWrapper_1_32 ZextWrapper_1_32_inst21(
    .I(ZextWrapper_1_32_inst21__I),
    .O(ZextWrapper_1_32_inst21__O)
  );

  wire [0:0] ZextWrapper_1_32_inst22__I;
  wire [31:0] ZextWrapper_1_32_inst22__O;
  ZextWrapper_1_32 ZextWrapper_1_32_inst22(
    .I(ZextWrapper_1_32_inst22__I),
    .O(ZextWrapper_1_32_inst22__O)
  );

  wire [0:0] ZextWrapper_1_32_inst23__I;
  wire [31:0] ZextWrapper_1_32_inst23__O;
  ZextWrapper_1_32 ZextWrapper_1_32_inst23(
    .I(ZextWrapper_1_32_inst23__I),
    .O(ZextWrapper_1_32_inst23__O)
  );

  wire [0:0] ZextWrapper_1_32_inst24__I;
  wire [31:0] ZextWrapper_1_32_inst24__O;
  ZextWrapper_1_32 ZextWrapper_1_32_inst24(
    .I(ZextWrapper_1_32_inst24__I),
    .O(ZextWrapper_1_32_inst24__O)
  );

  wire [0:0] ZextWrapper_1_32_inst25__I;
  wire [31:0] ZextWrapper_1_32_inst25__O;
  ZextWrapper_1_32 ZextWrapper_1_32_inst25(
    .I(ZextWrapper_1_32_inst25__I),
    .O(ZextWrapper_1_32_inst25__O)
  );

  wire [0:0] ZextWrapper_1_32_inst26__I;
  wire [31:0] ZextWrapper_1_32_inst26__O;
  ZextWrapper_1_32 ZextWrapper_1_32_inst26(
    .I(ZextWrapper_1_32_inst26__I),
    .O(ZextWrapper_1_32_inst26__O)
  );

  wire [0:0] ZextWrapper_1_32_inst27__I;
  wire [31:0] ZextWrapper_1_32_inst27__O;
  ZextWrapper_1_32 ZextWrapper_1_32_inst27(
    .I(ZextWrapper_1_32_inst27__I),
    .O(ZextWrapper_1_32_inst27__O)
  );

  wire [0:0] ZextWrapper_1_32_inst28__I;
  wire [31:0] ZextWrapper_1_32_inst28__O;
  ZextWrapper_1_32 ZextWrapper_1_32_inst28(
    .I(ZextWrapper_1_32_inst28__I),
    .O(ZextWrapper_1_32_inst28__O)
  );

  wire [0:0] ZextWrapper_1_32_inst29__I;
  wire [31:0] ZextWrapper_1_32_inst29__O;
  ZextWrapper_1_32 ZextWrapper_1_32_inst29(
    .I(ZextWrapper_1_32_inst29__I),
    .O(ZextWrapper_1_32_inst29__O)
  );

  wire [0:0] ZextWrapper_1_32_inst3__I;
  wire [31:0] ZextWrapper_1_32_inst3__O;
  ZextWrapper_1_32 ZextWrapper_1_32_inst3(
    .I(ZextWrapper_1_32_inst3__I),
    .O(ZextWrapper_1_32_inst3__O)
  );

  wire [0:0] ZextWrapper_1_32_inst30__I;
  wire [31:0] ZextWrapper_1_32_inst30__O;
  ZextWrapper_1_32 ZextWrapper_1_32_inst30(
    .I(ZextWrapper_1_32_inst30__I),
    .O(ZextWrapper_1_32_inst30__O)
  );

  wire [0:0] ZextWrapper_1_32_inst31__I;
  wire [31:0] ZextWrapper_1_32_inst31__O;
  ZextWrapper_1_32 ZextWrapper_1_32_inst31(
    .I(ZextWrapper_1_32_inst31__I),
    .O(ZextWrapper_1_32_inst31__O)
  );

  wire [0:0] ZextWrapper_1_32_inst32__I;
  wire [31:0] ZextWrapper_1_32_inst32__O;
  ZextWrapper_1_32 ZextWrapper_1_32_inst32(
    .I(ZextWrapper_1_32_inst32__I),
    .O(ZextWrapper_1_32_inst32__O)
  );

  wire [0:0] ZextWrapper_1_32_inst33__I;
  wire [31:0] ZextWrapper_1_32_inst33__O;
  ZextWrapper_1_32 ZextWrapper_1_32_inst33(
    .I(ZextWrapper_1_32_inst33__I),
    .O(ZextWrapper_1_32_inst33__O)
  );

  wire [0:0] ZextWrapper_1_32_inst34__I;
  wire [31:0] ZextWrapper_1_32_inst34__O;
  ZextWrapper_1_32 ZextWrapper_1_32_inst34(
    .I(ZextWrapper_1_32_inst34__I),
    .O(ZextWrapper_1_32_inst34__O)
  );

  wire [0:0] ZextWrapper_1_32_inst35__I;
  wire [31:0] ZextWrapper_1_32_inst35__O;
  ZextWrapper_1_32 ZextWrapper_1_32_inst35(
    .I(ZextWrapper_1_32_inst35__I),
    .O(ZextWrapper_1_32_inst35__O)
  );

  wire [0:0] ZextWrapper_1_32_inst36__I;
  wire [31:0] ZextWrapper_1_32_inst36__O;
  ZextWrapper_1_32 ZextWrapper_1_32_inst36(
    .I(ZextWrapper_1_32_inst36__I),
    .O(ZextWrapper_1_32_inst36__O)
  );

  wire [0:0] ZextWrapper_1_32_inst37__I;
  wire [31:0] ZextWrapper_1_32_inst37__O;
  ZextWrapper_1_32 ZextWrapper_1_32_inst37(
    .I(ZextWrapper_1_32_inst37__I),
    .O(ZextWrapper_1_32_inst37__O)
  );

  wire [0:0] ZextWrapper_1_32_inst38__I;
  wire [31:0] ZextWrapper_1_32_inst38__O;
  ZextWrapper_1_32 ZextWrapper_1_32_inst38(
    .I(ZextWrapper_1_32_inst38__I),
    .O(ZextWrapper_1_32_inst38__O)
  );

  wire [0:0] ZextWrapper_1_32_inst39__I;
  wire [31:0] ZextWrapper_1_32_inst39__O;
  ZextWrapper_1_32 ZextWrapper_1_32_inst39(
    .I(ZextWrapper_1_32_inst39__I),
    .O(ZextWrapper_1_32_inst39__O)
  );

  wire [0:0] ZextWrapper_1_32_inst4__I;
  wire [31:0] ZextWrapper_1_32_inst4__O;
  ZextWrapper_1_32 ZextWrapper_1_32_inst4(
    .I(ZextWrapper_1_32_inst4__I),
    .O(ZextWrapper_1_32_inst4__O)
  );

  wire [0:0] ZextWrapper_1_32_inst5__I;
  wire [31:0] ZextWrapper_1_32_inst5__O;
  ZextWrapper_1_32 ZextWrapper_1_32_inst5(
    .I(ZextWrapper_1_32_inst5__I),
    .O(ZextWrapper_1_32_inst5__O)
  );

  wire [0:0] ZextWrapper_1_32_inst6__I;
  wire [31:0] ZextWrapper_1_32_inst6__O;
  ZextWrapper_1_32 ZextWrapper_1_32_inst6(
    .I(ZextWrapper_1_32_inst6__I),
    .O(ZextWrapper_1_32_inst6__O)
  );

  wire [0:0] ZextWrapper_1_32_inst7__I;
  wire [31:0] ZextWrapper_1_32_inst7__O;
  ZextWrapper_1_32 ZextWrapper_1_32_inst7(
    .I(ZextWrapper_1_32_inst7__I),
    .O(ZextWrapper_1_32_inst7__O)
  );

  wire [0:0] ZextWrapper_1_32_inst8__I;
  wire [31:0] ZextWrapper_1_32_inst8__O;
  ZextWrapper_1_32 ZextWrapper_1_32_inst8(
    .I(ZextWrapper_1_32_inst8__I),
    .O(ZextWrapper_1_32_inst8__O)
  );

  wire [0:0] ZextWrapper_1_32_inst9__I;
  wire [31:0] ZextWrapper_1_32_inst9__O;
  ZextWrapper_1_32 ZextWrapper_1_32_inst9(
    .I(ZextWrapper_1_32_inst9__I),
    .O(ZextWrapper_1_32_inst9__O)
  );

  wire [1:0] ZextWrapper_2_32_inst0__I;
  wire [31:0] ZextWrapper_2_32_inst0__O;
  ZextWrapper_2_32 ZextWrapper_2_32_inst0(
    .I(ZextWrapper_2_32_inst0__I),
    .O(ZextWrapper_2_32_inst0__O)
  );

  wire [1:0] ZextWrapper_2_32_inst1__I;
  wire [31:0] ZextWrapper_2_32_inst1__O;
  ZextWrapper_2_32 ZextWrapper_2_32_inst1(
    .I(ZextWrapper_2_32_inst1__I),
    .O(ZextWrapper_2_32_inst1__O)
  );

  wire [1:0] ZextWrapper_2_32_inst10__I;
  wire [31:0] ZextWrapper_2_32_inst10__O;
  ZextWrapper_2_32 ZextWrapper_2_32_inst10(
    .I(ZextWrapper_2_32_inst10__I),
    .O(ZextWrapper_2_32_inst10__O)
  );

  wire [1:0] ZextWrapper_2_32_inst11__I;
  wire [31:0] ZextWrapper_2_32_inst11__O;
  ZextWrapper_2_32 ZextWrapper_2_32_inst11(
    .I(ZextWrapper_2_32_inst11__I),
    .O(ZextWrapper_2_32_inst11__O)
  );

  wire [1:0] ZextWrapper_2_32_inst12__I;
  wire [31:0] ZextWrapper_2_32_inst12__O;
  ZextWrapper_2_32 ZextWrapper_2_32_inst12(
    .I(ZextWrapper_2_32_inst12__I),
    .O(ZextWrapper_2_32_inst12__O)
  );

  wire [1:0] ZextWrapper_2_32_inst13__I;
  wire [31:0] ZextWrapper_2_32_inst13__O;
  ZextWrapper_2_32 ZextWrapper_2_32_inst13(
    .I(ZextWrapper_2_32_inst13__I),
    .O(ZextWrapper_2_32_inst13__O)
  );

  wire [1:0] ZextWrapper_2_32_inst14__I;
  wire [31:0] ZextWrapper_2_32_inst14__O;
  ZextWrapper_2_32 ZextWrapper_2_32_inst14(
    .I(ZextWrapper_2_32_inst14__I),
    .O(ZextWrapper_2_32_inst14__O)
  );

  wire [1:0] ZextWrapper_2_32_inst15__I;
  wire [31:0] ZextWrapper_2_32_inst15__O;
  ZextWrapper_2_32 ZextWrapper_2_32_inst15(
    .I(ZextWrapper_2_32_inst15__I),
    .O(ZextWrapper_2_32_inst15__O)
  );

  wire [1:0] ZextWrapper_2_32_inst16__I;
  wire [31:0] ZextWrapper_2_32_inst16__O;
  ZextWrapper_2_32 ZextWrapper_2_32_inst16(
    .I(ZextWrapper_2_32_inst16__I),
    .O(ZextWrapper_2_32_inst16__O)
  );

  wire [1:0] ZextWrapper_2_32_inst17__I;
  wire [31:0] ZextWrapper_2_32_inst17__O;
  ZextWrapper_2_32 ZextWrapper_2_32_inst17(
    .I(ZextWrapper_2_32_inst17__I),
    .O(ZextWrapper_2_32_inst17__O)
  );

  wire [1:0] ZextWrapper_2_32_inst18__I;
  wire [31:0] ZextWrapper_2_32_inst18__O;
  ZextWrapper_2_32 ZextWrapper_2_32_inst18(
    .I(ZextWrapper_2_32_inst18__I),
    .O(ZextWrapper_2_32_inst18__O)
  );

  wire [1:0] ZextWrapper_2_32_inst19__I;
  wire [31:0] ZextWrapper_2_32_inst19__O;
  ZextWrapper_2_32 ZextWrapper_2_32_inst19(
    .I(ZextWrapper_2_32_inst19__I),
    .O(ZextWrapper_2_32_inst19__O)
  );

  wire [1:0] ZextWrapper_2_32_inst2__I;
  wire [31:0] ZextWrapper_2_32_inst2__O;
  ZextWrapper_2_32 ZextWrapper_2_32_inst2(
    .I(ZextWrapper_2_32_inst2__I),
    .O(ZextWrapper_2_32_inst2__O)
  );

  wire [1:0] ZextWrapper_2_32_inst20__I;
  wire [31:0] ZextWrapper_2_32_inst20__O;
  ZextWrapper_2_32 ZextWrapper_2_32_inst20(
    .I(ZextWrapper_2_32_inst20__I),
    .O(ZextWrapper_2_32_inst20__O)
  );

  wire [1:0] ZextWrapper_2_32_inst21__I;
  wire [31:0] ZextWrapper_2_32_inst21__O;
  ZextWrapper_2_32 ZextWrapper_2_32_inst21(
    .I(ZextWrapper_2_32_inst21__I),
    .O(ZextWrapper_2_32_inst21__O)
  );

  wire [1:0] ZextWrapper_2_32_inst22__I;
  wire [31:0] ZextWrapper_2_32_inst22__O;
  ZextWrapper_2_32 ZextWrapper_2_32_inst22(
    .I(ZextWrapper_2_32_inst22__I),
    .O(ZextWrapper_2_32_inst22__O)
  );

  wire [1:0] ZextWrapper_2_32_inst23__I;
  wire [31:0] ZextWrapper_2_32_inst23__O;
  ZextWrapper_2_32 ZextWrapper_2_32_inst23(
    .I(ZextWrapper_2_32_inst23__I),
    .O(ZextWrapper_2_32_inst23__O)
  );

  wire [1:0] ZextWrapper_2_32_inst24__I;
  wire [31:0] ZextWrapper_2_32_inst24__O;
  ZextWrapper_2_32 ZextWrapper_2_32_inst24(
    .I(ZextWrapper_2_32_inst24__I),
    .O(ZextWrapper_2_32_inst24__O)
  );

  wire [1:0] ZextWrapper_2_32_inst25__I;
  wire [31:0] ZextWrapper_2_32_inst25__O;
  ZextWrapper_2_32 ZextWrapper_2_32_inst25(
    .I(ZextWrapper_2_32_inst25__I),
    .O(ZextWrapper_2_32_inst25__O)
  );

  wire [1:0] ZextWrapper_2_32_inst26__I;
  wire [31:0] ZextWrapper_2_32_inst26__O;
  ZextWrapper_2_32 ZextWrapper_2_32_inst26(
    .I(ZextWrapper_2_32_inst26__I),
    .O(ZextWrapper_2_32_inst26__O)
  );

  wire [1:0] ZextWrapper_2_32_inst27__I;
  wire [31:0] ZextWrapper_2_32_inst27__O;
  ZextWrapper_2_32 ZextWrapper_2_32_inst27(
    .I(ZextWrapper_2_32_inst27__I),
    .O(ZextWrapper_2_32_inst27__O)
  );

  wire [1:0] ZextWrapper_2_32_inst28__I;
  wire [31:0] ZextWrapper_2_32_inst28__O;
  ZextWrapper_2_32 ZextWrapper_2_32_inst28(
    .I(ZextWrapper_2_32_inst28__I),
    .O(ZextWrapper_2_32_inst28__O)
  );

  wire [1:0] ZextWrapper_2_32_inst29__I;
  wire [31:0] ZextWrapper_2_32_inst29__O;
  ZextWrapper_2_32 ZextWrapper_2_32_inst29(
    .I(ZextWrapper_2_32_inst29__I),
    .O(ZextWrapper_2_32_inst29__O)
  );

  wire [1:0] ZextWrapper_2_32_inst3__I;
  wire [31:0] ZextWrapper_2_32_inst3__O;
  ZextWrapper_2_32 ZextWrapper_2_32_inst3(
    .I(ZextWrapper_2_32_inst3__I),
    .O(ZextWrapper_2_32_inst3__O)
  );

  wire [1:0] ZextWrapper_2_32_inst30__I;
  wire [31:0] ZextWrapper_2_32_inst30__O;
  ZextWrapper_2_32 ZextWrapper_2_32_inst30(
    .I(ZextWrapper_2_32_inst30__I),
    .O(ZextWrapper_2_32_inst30__O)
  );

  wire [1:0] ZextWrapper_2_32_inst31__I;
  wire [31:0] ZextWrapper_2_32_inst31__O;
  ZextWrapper_2_32 ZextWrapper_2_32_inst31(
    .I(ZextWrapper_2_32_inst31__I),
    .O(ZextWrapper_2_32_inst31__O)
  );

  wire [1:0] ZextWrapper_2_32_inst32__I;
  wire [31:0] ZextWrapper_2_32_inst32__O;
  ZextWrapper_2_32 ZextWrapper_2_32_inst32(
    .I(ZextWrapper_2_32_inst32__I),
    .O(ZextWrapper_2_32_inst32__O)
  );

  wire [1:0] ZextWrapper_2_32_inst33__I;
  wire [31:0] ZextWrapper_2_32_inst33__O;
  ZextWrapper_2_32 ZextWrapper_2_32_inst33(
    .I(ZextWrapper_2_32_inst33__I),
    .O(ZextWrapper_2_32_inst33__O)
  );

  wire [1:0] ZextWrapper_2_32_inst34__I;
  wire [31:0] ZextWrapper_2_32_inst34__O;
  ZextWrapper_2_32 ZextWrapper_2_32_inst34(
    .I(ZextWrapper_2_32_inst34__I),
    .O(ZextWrapper_2_32_inst34__O)
  );

  wire [1:0] ZextWrapper_2_32_inst35__I;
  wire [31:0] ZextWrapper_2_32_inst35__O;
  ZextWrapper_2_32 ZextWrapper_2_32_inst35(
    .I(ZextWrapper_2_32_inst35__I),
    .O(ZextWrapper_2_32_inst35__O)
  );

  wire [1:0] ZextWrapper_2_32_inst36__I;
  wire [31:0] ZextWrapper_2_32_inst36__O;
  ZextWrapper_2_32 ZextWrapper_2_32_inst36(
    .I(ZextWrapper_2_32_inst36__I),
    .O(ZextWrapper_2_32_inst36__O)
  );

  wire [1:0] ZextWrapper_2_32_inst37__I;
  wire [31:0] ZextWrapper_2_32_inst37__O;
  ZextWrapper_2_32 ZextWrapper_2_32_inst37(
    .I(ZextWrapper_2_32_inst37__I),
    .O(ZextWrapper_2_32_inst37__O)
  );

  wire [1:0] ZextWrapper_2_32_inst38__I;
  wire [31:0] ZextWrapper_2_32_inst38__O;
  ZextWrapper_2_32 ZextWrapper_2_32_inst38(
    .I(ZextWrapper_2_32_inst38__I),
    .O(ZextWrapper_2_32_inst38__O)
  );

  wire [1:0] ZextWrapper_2_32_inst39__I;
  wire [31:0] ZextWrapper_2_32_inst39__O;
  ZextWrapper_2_32 ZextWrapper_2_32_inst39(
    .I(ZextWrapper_2_32_inst39__I),
    .O(ZextWrapper_2_32_inst39__O)
  );

  wire [1:0] ZextWrapper_2_32_inst4__I;
  wire [31:0] ZextWrapper_2_32_inst4__O;
  ZextWrapper_2_32 ZextWrapper_2_32_inst4(
    .I(ZextWrapper_2_32_inst4__I),
    .O(ZextWrapper_2_32_inst4__O)
  );

  wire [1:0] ZextWrapper_2_32_inst5__I;
  wire [31:0] ZextWrapper_2_32_inst5__O;
  ZextWrapper_2_32 ZextWrapper_2_32_inst5(
    .I(ZextWrapper_2_32_inst5__I),
    .O(ZextWrapper_2_32_inst5__O)
  );

  wire [1:0] ZextWrapper_2_32_inst6__I;
  wire [31:0] ZextWrapper_2_32_inst6__O;
  ZextWrapper_2_32 ZextWrapper_2_32_inst6(
    .I(ZextWrapper_2_32_inst6__I),
    .O(ZextWrapper_2_32_inst6__O)
  );

  wire [1:0] ZextWrapper_2_32_inst7__I;
  wire [31:0] ZextWrapper_2_32_inst7__O;
  ZextWrapper_2_32 ZextWrapper_2_32_inst7(
    .I(ZextWrapper_2_32_inst7__I),
    .O(ZextWrapper_2_32_inst7__O)
  );

  wire [1:0] ZextWrapper_2_32_inst8__I;
  wire [31:0] ZextWrapper_2_32_inst8__O;
  ZextWrapper_2_32 ZextWrapper_2_32_inst8(
    .I(ZextWrapper_2_32_inst8__I),
    .O(ZextWrapper_2_32_inst8__O)
  );

  wire [1:0] ZextWrapper_2_32_inst9__I;
  wire [31:0] ZextWrapper_2_32_inst9__O;
  ZextWrapper_2_32 ZextWrapper_2_32_inst9(
    .I(ZextWrapper_2_32_inst9__I),
    .O(ZextWrapper_2_32_inst9__O)
  );

  // Instancing generated Module: coreir.reg(width:1)
  wire  reg_P_inst0__clk;
  wire [0:0] reg_P_inst0__in;
  wire [0:0] reg_P_inst0__out;
  coreir_reg #(.clk_posedge(1),.init(1'h0),.width(1)) reg_P_inst0(
    .clk(reg_P_inst0__clk),
    .in(reg_P_inst0__in),
    .out(reg_P_inst0__out)
  );

  // Instancing generated Module: coreir.reg(width:1)
  wire  reg_P_inst1__clk;
  wire [0:0] reg_P_inst1__in;
  wire [0:0] reg_P_inst1__out;
  coreir_reg #(.clk_posedge(1),.init(1'h0),.width(1)) reg_P_inst1(
    .clk(reg_P_inst1__clk),
    .in(reg_P_inst1__in),
    .out(reg_P_inst1__out)
  );

  // Instancing generated Module: coreir.reg(width:1)
  wire  reg_P_inst10__clk;
  wire [0:0] reg_P_inst10__in;
  wire [0:0] reg_P_inst10__out;
  coreir_reg #(.clk_posedge(1),.init(1'h0),.width(1)) reg_P_inst10(
    .clk(reg_P_inst10__clk),
    .in(reg_P_inst10__in),
    .out(reg_P_inst10__out)
  );

  // Instancing generated Module: coreir.reg(width:1)
  wire  reg_P_inst11__clk;
  wire [0:0] reg_P_inst11__in;
  wire [0:0] reg_P_inst11__out;
  coreir_reg #(.clk_posedge(1),.init(1'h0),.width(1)) reg_P_inst11(
    .clk(reg_P_inst11__clk),
    .in(reg_P_inst11__in),
    .out(reg_P_inst11__out)
  );

  // Instancing generated Module: coreir.reg(width:1)
  wire  reg_P_inst12__clk;
  wire [0:0] reg_P_inst12__in;
  wire [0:0] reg_P_inst12__out;
  coreir_reg #(.clk_posedge(1),.init(1'h0),.width(1)) reg_P_inst12(
    .clk(reg_P_inst12__clk),
    .in(reg_P_inst12__in),
    .out(reg_P_inst12__out)
  );

  // Instancing generated Module: coreir.reg(width:1)
  wire  reg_P_inst13__clk;
  wire [0:0] reg_P_inst13__in;
  wire [0:0] reg_P_inst13__out;
  coreir_reg #(.clk_posedge(1),.init(1'h0),.width(1)) reg_P_inst13(
    .clk(reg_P_inst13__clk),
    .in(reg_P_inst13__in),
    .out(reg_P_inst13__out)
  );

  // Instancing generated Module: coreir.reg(width:1)
  wire  reg_P_inst14__clk;
  wire [0:0] reg_P_inst14__in;
  wire [0:0] reg_P_inst14__out;
  coreir_reg #(.clk_posedge(1),.init(1'h0),.width(1)) reg_P_inst14(
    .clk(reg_P_inst14__clk),
    .in(reg_P_inst14__in),
    .out(reg_P_inst14__out)
  );

  // Instancing generated Module: coreir.reg(width:16)
  wire  reg_P_inst15__clk;
  wire [15:0] reg_P_inst15__in;
  wire [15:0] reg_P_inst15__out;
  coreir_reg #(.clk_posedge(1),.init(16'h0000),.width(16)) reg_P_inst15(
    .clk(reg_P_inst15__clk),
    .in(reg_P_inst15__in),
    .out(reg_P_inst15__out)
  );

  // Instancing generated Module: coreir.reg(width:16)
  wire  reg_P_inst16__clk;
  wire [15:0] reg_P_inst16__in;
  wire [15:0] reg_P_inst16__out;
  coreir_reg #(.clk_posedge(1),.init(16'h0000),.width(16)) reg_P_inst16(
    .clk(reg_P_inst16__clk),
    .in(reg_P_inst16__in),
    .out(reg_P_inst16__out)
  );

  // Instancing generated Module: coreir.reg(width:16)
  wire  reg_P_inst17__clk;
  wire [15:0] reg_P_inst17__in;
  wire [15:0] reg_P_inst17__out;
  coreir_reg #(.clk_posedge(1),.init(16'h0000),.width(16)) reg_P_inst17(
    .clk(reg_P_inst17__clk),
    .in(reg_P_inst17__in),
    .out(reg_P_inst17__out)
  );

  // Instancing generated Module: coreir.reg(width:16)
  wire  reg_P_inst18__clk;
  wire [15:0] reg_P_inst18__in;
  wire [15:0] reg_P_inst18__out;
  coreir_reg #(.clk_posedge(1),.init(16'h0000),.width(16)) reg_P_inst18(
    .clk(reg_P_inst18__clk),
    .in(reg_P_inst18__in),
    .out(reg_P_inst18__out)
  );

  // Instancing generated Module: coreir.reg(width:16)
  wire  reg_P_inst19__clk;
  wire [15:0] reg_P_inst19__in;
  wire [15:0] reg_P_inst19__out;
  coreir_reg #(.clk_posedge(1),.init(16'h0000),.width(16)) reg_P_inst19(
    .clk(reg_P_inst19__clk),
    .in(reg_P_inst19__in),
    .out(reg_P_inst19__out)
  );

  // Instancing generated Module: coreir.reg(width:1)
  wire  reg_P_inst2__clk;
  wire [0:0] reg_P_inst2__in;
  wire [0:0] reg_P_inst2__out;
  coreir_reg #(.clk_posedge(1),.init(1'h0),.width(1)) reg_P_inst2(
    .clk(reg_P_inst2__clk),
    .in(reg_P_inst2__in),
    .out(reg_P_inst2__out)
  );

  // Instancing generated Module: coreir.reg(width:1)
  wire  reg_P_inst20__clk;
  wire [0:0] reg_P_inst20__in;
  wire [0:0] reg_P_inst20__out;
  coreir_reg #(.clk_posedge(1),.init(1'h0),.width(1)) reg_P_inst20(
    .clk(reg_P_inst20__clk),
    .in(reg_P_inst20__in),
    .out(reg_P_inst20__out)
  );

  // Instancing generated Module: coreir.reg(width:1)
  wire  reg_P_inst21__clk;
  wire [0:0] reg_P_inst21__in;
  wire [0:0] reg_P_inst21__out;
  coreir_reg #(.clk_posedge(1),.init(1'h0),.width(1)) reg_P_inst21(
    .clk(reg_P_inst21__clk),
    .in(reg_P_inst21__in),
    .out(reg_P_inst21__out)
  );

  // Instancing generated Module: coreir.reg(width:1)
  wire  reg_P_inst22__clk;
  wire [0:0] reg_P_inst22__in;
  wire [0:0] reg_P_inst22__out;
  coreir_reg #(.clk_posedge(1),.init(1'h0),.width(1)) reg_P_inst22(
    .clk(reg_P_inst22__clk),
    .in(reg_P_inst22__in),
    .out(reg_P_inst22__out)
  );

  // Instancing generated Module: coreir.reg(width:1)
  wire  reg_P_inst23__clk;
  wire [0:0] reg_P_inst23__in;
  wire [0:0] reg_P_inst23__out;
  coreir_reg #(.clk_posedge(1),.init(1'h0),.width(1)) reg_P_inst23(
    .clk(reg_P_inst23__clk),
    .in(reg_P_inst23__in),
    .out(reg_P_inst23__out)
  );

  // Instancing generated Module: coreir.reg(width:1)
  wire  reg_P_inst24__clk;
  wire [0:0] reg_P_inst24__in;
  wire [0:0] reg_P_inst24__out;
  coreir_reg #(.clk_posedge(1),.init(1'h0),.width(1)) reg_P_inst24(
    .clk(reg_P_inst24__clk),
    .in(reg_P_inst24__in),
    .out(reg_P_inst24__out)
  );

  // Instancing generated Module: coreir.reg(width:16)
  wire  reg_P_inst25__clk;
  wire [15:0] reg_P_inst25__in;
  wire [15:0] reg_P_inst25__out;
  coreir_reg #(.clk_posedge(1),.init(16'h0000),.width(16)) reg_P_inst25(
    .clk(reg_P_inst25__clk),
    .in(reg_P_inst25__in),
    .out(reg_P_inst25__out)
  );

  // Instancing generated Module: coreir.reg(width:16)
  wire  reg_P_inst26__clk;
  wire [15:0] reg_P_inst26__in;
  wire [15:0] reg_P_inst26__out;
  coreir_reg #(.clk_posedge(1),.init(16'h0000),.width(16)) reg_P_inst26(
    .clk(reg_P_inst26__clk),
    .in(reg_P_inst26__in),
    .out(reg_P_inst26__out)
  );

  // Instancing generated Module: coreir.reg(width:16)
  wire  reg_P_inst27__clk;
  wire [15:0] reg_P_inst27__in;
  wire [15:0] reg_P_inst27__out;
  coreir_reg #(.clk_posedge(1),.init(16'h0000),.width(16)) reg_P_inst27(
    .clk(reg_P_inst27__clk),
    .in(reg_P_inst27__in),
    .out(reg_P_inst27__out)
  );

  // Instancing generated Module: coreir.reg(width:16)
  wire  reg_P_inst28__clk;
  wire [15:0] reg_P_inst28__in;
  wire [15:0] reg_P_inst28__out;
  coreir_reg #(.clk_posedge(1),.init(16'h0000),.width(16)) reg_P_inst28(
    .clk(reg_P_inst28__clk),
    .in(reg_P_inst28__in),
    .out(reg_P_inst28__out)
  );

  // Instancing generated Module: coreir.reg(width:16)
  wire  reg_P_inst29__clk;
  wire [15:0] reg_P_inst29__in;
  wire [15:0] reg_P_inst29__out;
  coreir_reg #(.clk_posedge(1),.init(16'h0000),.width(16)) reg_P_inst29(
    .clk(reg_P_inst29__clk),
    .in(reg_P_inst29__in),
    .out(reg_P_inst29__out)
  );

  // Instancing generated Module: coreir.reg(width:1)
  wire  reg_P_inst3__clk;
  wire [0:0] reg_P_inst3__in;
  wire [0:0] reg_P_inst3__out;
  coreir_reg #(.clk_posedge(1),.init(1'h0),.width(1)) reg_P_inst3(
    .clk(reg_P_inst3__clk),
    .in(reg_P_inst3__in),
    .out(reg_P_inst3__out)
  );

  // Instancing generated Module: coreir.reg(width:1)
  wire  reg_P_inst30__clk;
  wire [0:0] reg_P_inst30__in;
  wire [0:0] reg_P_inst30__out;
  coreir_reg #(.clk_posedge(1),.init(1'h0),.width(1)) reg_P_inst30(
    .clk(reg_P_inst30__clk),
    .in(reg_P_inst30__in),
    .out(reg_P_inst30__out)
  );

  // Instancing generated Module: coreir.reg(width:1)
  wire  reg_P_inst31__clk;
  wire [0:0] reg_P_inst31__in;
  wire [0:0] reg_P_inst31__out;
  coreir_reg #(.clk_posedge(1),.init(1'h0),.width(1)) reg_P_inst31(
    .clk(reg_P_inst31__clk),
    .in(reg_P_inst31__in),
    .out(reg_P_inst31__out)
  );

  // Instancing generated Module: coreir.reg(width:1)
  wire  reg_P_inst32__clk;
  wire [0:0] reg_P_inst32__in;
  wire [0:0] reg_P_inst32__out;
  coreir_reg #(.clk_posedge(1),.init(1'h0),.width(1)) reg_P_inst32(
    .clk(reg_P_inst32__clk),
    .in(reg_P_inst32__in),
    .out(reg_P_inst32__out)
  );

  // Instancing generated Module: coreir.reg(width:1)
  wire  reg_P_inst33__clk;
  wire [0:0] reg_P_inst33__in;
  wire [0:0] reg_P_inst33__out;
  coreir_reg #(.clk_posedge(1),.init(1'h0),.width(1)) reg_P_inst33(
    .clk(reg_P_inst33__clk),
    .in(reg_P_inst33__in),
    .out(reg_P_inst33__out)
  );

  // Instancing generated Module: coreir.reg(width:1)
  wire  reg_P_inst34__clk;
  wire [0:0] reg_P_inst34__in;
  wire [0:0] reg_P_inst34__out;
  coreir_reg #(.clk_posedge(1),.init(1'h0),.width(1)) reg_P_inst34(
    .clk(reg_P_inst34__clk),
    .in(reg_P_inst34__in),
    .out(reg_P_inst34__out)
  );

  // Instancing generated Module: coreir.reg(width:16)
  wire  reg_P_inst35__clk;
  wire [15:0] reg_P_inst35__in;
  wire [15:0] reg_P_inst35__out;
  coreir_reg #(.clk_posedge(1),.init(16'h0000),.width(16)) reg_P_inst35(
    .clk(reg_P_inst35__clk),
    .in(reg_P_inst35__in),
    .out(reg_P_inst35__out)
  );

  // Instancing generated Module: coreir.reg(width:16)
  wire  reg_P_inst36__clk;
  wire [15:0] reg_P_inst36__in;
  wire [15:0] reg_P_inst36__out;
  coreir_reg #(.clk_posedge(1),.init(16'h0000),.width(16)) reg_P_inst36(
    .clk(reg_P_inst36__clk),
    .in(reg_P_inst36__in),
    .out(reg_P_inst36__out)
  );

  // Instancing generated Module: coreir.reg(width:16)
  wire  reg_P_inst37__clk;
  wire [15:0] reg_P_inst37__in;
  wire [15:0] reg_P_inst37__out;
  coreir_reg #(.clk_posedge(1),.init(16'h0000),.width(16)) reg_P_inst37(
    .clk(reg_P_inst37__clk),
    .in(reg_P_inst37__in),
    .out(reg_P_inst37__out)
  );

  // Instancing generated Module: coreir.reg(width:16)
  wire  reg_P_inst38__clk;
  wire [15:0] reg_P_inst38__in;
  wire [15:0] reg_P_inst38__out;
  coreir_reg #(.clk_posedge(1),.init(16'h0000),.width(16)) reg_P_inst38(
    .clk(reg_P_inst38__clk),
    .in(reg_P_inst38__in),
    .out(reg_P_inst38__out)
  );

  // Instancing generated Module: coreir.reg(width:16)
  wire  reg_P_inst39__clk;
  wire [15:0] reg_P_inst39__in;
  wire [15:0] reg_P_inst39__out;
  coreir_reg #(.clk_posedge(1),.init(16'h0000),.width(16)) reg_P_inst39(
    .clk(reg_P_inst39__clk),
    .in(reg_P_inst39__in),
    .out(reg_P_inst39__out)
  );

  // Instancing generated Module: coreir.reg(width:1)
  wire  reg_P_inst4__clk;
  wire [0:0] reg_P_inst4__in;
  wire [0:0] reg_P_inst4__out;
  coreir_reg #(.clk_posedge(1),.init(1'h0),.width(1)) reg_P_inst4(
    .clk(reg_P_inst4__clk),
    .in(reg_P_inst4__in),
    .out(reg_P_inst4__out)
  );

  // Instancing generated Module: coreir.reg(width:16)
  wire  reg_P_inst5__clk;
  wire [15:0] reg_P_inst5__in;
  wire [15:0] reg_P_inst5__out;
  coreir_reg #(.clk_posedge(1),.init(16'h0000),.width(16)) reg_P_inst5(
    .clk(reg_P_inst5__clk),
    .in(reg_P_inst5__in),
    .out(reg_P_inst5__out)
  );

  // Instancing generated Module: coreir.reg(width:16)
  wire  reg_P_inst6__clk;
  wire [15:0] reg_P_inst6__in;
  wire [15:0] reg_P_inst6__out;
  coreir_reg #(.clk_posedge(1),.init(16'h0000),.width(16)) reg_P_inst6(
    .clk(reg_P_inst6__clk),
    .in(reg_P_inst6__in),
    .out(reg_P_inst6__out)
  );

  // Instancing generated Module: coreir.reg(width:16)
  wire  reg_P_inst7__clk;
  wire [15:0] reg_P_inst7__in;
  wire [15:0] reg_P_inst7__out;
  coreir_reg #(.clk_posedge(1),.init(16'h0000),.width(16)) reg_P_inst7(
    .clk(reg_P_inst7__clk),
    .in(reg_P_inst7__in),
    .out(reg_P_inst7__out)
  );

  // Instancing generated Module: coreir.reg(width:16)
  wire  reg_P_inst8__clk;
  wire [15:0] reg_P_inst8__in;
  wire [15:0] reg_P_inst8__out;
  coreir_reg #(.clk_posedge(1),.init(16'h0000),.width(16)) reg_P_inst8(
    .clk(reg_P_inst8__clk),
    .in(reg_P_inst8__in),
    .out(reg_P_inst8__out)
  );

  // Instancing generated Module: coreir.reg(width:16)
  wire  reg_P_inst9__clk;
  wire [15:0] reg_P_inst9__in;
  wire [15:0] reg_P_inst9__out;
  coreir_reg #(.clk_posedge(1),.init(16'h0000),.width(16)) reg_P_inst9(
    .clk(reg_P_inst9__clk),
    .in(reg_P_inst9__in),
    .out(reg_P_inst9__out)
  );

  assign MuxWrapper_2_16_inst0__S[0:0] = ConfigRegister_1_8_32_11_inst0__O[0:0];

  assign ZextWrapper_1_32_inst5__I[0:0] = ConfigRegister_1_8_32_11_inst0__O[0:0];

  assign ConfigRegister_1_8_32_11_inst0__clk = clk;

  assign ConfigRegister_1_8_32_11_inst0__config_addr[7:0] = config_config_addr[7:0];

  assign ConfigRegister_1_8_32_11_inst0__config_data[31:0] = config_config_data[31:0];

  assign ConfigRegister_1_8_32_11_inst0__config_en = config_write[0];

  assign ConfigRegister_1_8_32_11_inst0__reset = reset;

  assign MuxWrapper_2_16_inst1__S[0:0] = ConfigRegister_1_8_32_13_inst0__O[0:0];

  assign ZextWrapper_1_32_inst6__I[0:0] = ConfigRegister_1_8_32_13_inst0__O[0:0];

  assign ConfigRegister_1_8_32_13_inst0__clk = clk;

  assign ConfigRegister_1_8_32_13_inst0__config_addr[7:0] = config_config_addr[7:0];

  assign ConfigRegister_1_8_32_13_inst0__config_data[31:0] = config_config_data[31:0];

  assign ConfigRegister_1_8_32_13_inst0__config_en = config_write[0];

  assign ConfigRegister_1_8_32_13_inst0__reset = reset;

  assign MuxWrapper_2_16_inst2__S[0:0] = ConfigRegister_1_8_32_15_inst0__O[0:0];

  assign ZextWrapper_1_32_inst7__I[0:0] = ConfigRegister_1_8_32_15_inst0__O[0:0];

  assign ConfigRegister_1_8_32_15_inst0__clk = clk;

  assign ConfigRegister_1_8_32_15_inst0__config_addr[7:0] = config_config_addr[7:0];

  assign ConfigRegister_1_8_32_15_inst0__config_data[31:0] = config_config_data[31:0];

  assign ConfigRegister_1_8_32_15_inst0__config_en = config_write[0];

  assign ConfigRegister_1_8_32_15_inst0__reset = reset;

  assign MuxWrapper_2_16_inst3__S[0:0] = ConfigRegister_1_8_32_17_inst0__O[0:0];

  assign ZextWrapper_1_32_inst8__I[0:0] = ConfigRegister_1_8_32_17_inst0__O[0:0];

  assign ConfigRegister_1_8_32_17_inst0__clk = clk;

  assign ConfigRegister_1_8_32_17_inst0__config_addr[7:0] = config_config_addr[7:0];

  assign ConfigRegister_1_8_32_17_inst0__config_data[31:0] = config_config_data[31:0];

  assign ConfigRegister_1_8_32_17_inst0__config_en = config_write[0];

  assign ConfigRegister_1_8_32_17_inst0__reset = reset;

  assign MuxWrapper_2_16_inst4__S[0:0] = ConfigRegister_1_8_32_19_inst0__O[0:0];

  assign ZextWrapper_1_32_inst9__I[0:0] = ConfigRegister_1_8_32_19_inst0__O[0:0];

  assign ConfigRegister_1_8_32_19_inst0__clk = clk;

  assign ConfigRegister_1_8_32_19_inst0__config_addr[7:0] = config_config_addr[7:0];

  assign ConfigRegister_1_8_32_19_inst0__config_data[31:0] = config_config_data[31:0];

  assign ConfigRegister_1_8_32_19_inst0__config_en = config_write[0];

  assign ConfigRegister_1_8_32_19_inst0__reset = reset;

  assign MuxWrapper_2_1_inst0__S[0:0] = ConfigRegister_1_8_32_1_inst0__O[0:0];

  assign ZextWrapper_1_32_inst0__I[0:0] = ConfigRegister_1_8_32_1_inst0__O[0:0];

  assign ConfigRegister_1_8_32_1_inst0__clk = clk;

  assign ConfigRegister_1_8_32_1_inst0__config_addr[7:0] = config_config_addr[7:0];

  assign ConfigRegister_1_8_32_1_inst0__config_data[31:0] = config_config_data[31:0];

  assign ConfigRegister_1_8_32_1_inst0__config_en = config_write[0];

  assign ConfigRegister_1_8_32_1_inst0__reset = reset;

  assign MuxWrapper_2_1_inst5__S[0:0] = ConfigRegister_1_8_32_21_inst0__O[0:0];

  assign ZextWrapper_1_32_inst10__I[0:0] = ConfigRegister_1_8_32_21_inst0__O[0:0];

  assign ConfigRegister_1_8_32_21_inst0__clk = clk;

  assign ConfigRegister_1_8_32_21_inst0__config_addr[7:0] = config_config_addr[7:0];

  assign ConfigRegister_1_8_32_21_inst0__config_data[31:0] = config_config_data[31:0];

  assign ConfigRegister_1_8_32_21_inst0__config_en = config_write[0];

  assign ConfigRegister_1_8_32_21_inst0__reset = reset;

  assign MuxWrapper_2_1_inst6__S[0:0] = ConfigRegister_1_8_32_23_inst0__O[0:0];

  assign ZextWrapper_1_32_inst11__I[0:0] = ConfigRegister_1_8_32_23_inst0__O[0:0];

  assign ConfigRegister_1_8_32_23_inst0__clk = clk;

  assign ConfigRegister_1_8_32_23_inst0__config_addr[7:0] = config_config_addr[7:0];

  assign ConfigRegister_1_8_32_23_inst0__config_data[31:0] = config_config_data[31:0];

  assign ConfigRegister_1_8_32_23_inst0__config_en = config_write[0];

  assign ConfigRegister_1_8_32_23_inst0__reset = reset;

  assign MuxWrapper_2_1_inst7__S[0:0] = ConfigRegister_1_8_32_25_inst0__O[0:0];

  assign ZextWrapper_1_32_inst12__I[0:0] = ConfigRegister_1_8_32_25_inst0__O[0:0];

  assign ConfigRegister_1_8_32_25_inst0__clk = clk;

  assign ConfigRegister_1_8_32_25_inst0__config_addr[7:0] = config_config_addr[7:0];

  assign ConfigRegister_1_8_32_25_inst0__config_data[31:0] = config_config_data[31:0];

  assign ConfigRegister_1_8_32_25_inst0__config_en = config_write[0];

  assign ConfigRegister_1_8_32_25_inst0__reset = reset;

  assign MuxWrapper_2_1_inst8__S[0:0] = ConfigRegister_1_8_32_27_inst0__O[0:0];

  assign ZextWrapper_1_32_inst13__I[0:0] = ConfigRegister_1_8_32_27_inst0__O[0:0];

  assign ConfigRegister_1_8_32_27_inst0__clk = clk;

  assign ConfigRegister_1_8_32_27_inst0__config_addr[7:0] = config_config_addr[7:0];

  assign ConfigRegister_1_8_32_27_inst0__config_data[31:0] = config_config_data[31:0];

  assign ConfigRegister_1_8_32_27_inst0__config_en = config_write[0];

  assign ConfigRegister_1_8_32_27_inst0__reset = reset;

  assign MuxWrapper_2_1_inst9__S[0:0] = ConfigRegister_1_8_32_29_inst0__O[0:0];

  assign ZextWrapper_1_32_inst14__I[0:0] = ConfigRegister_1_8_32_29_inst0__O[0:0];

  assign ConfigRegister_1_8_32_29_inst0__clk = clk;

  assign ConfigRegister_1_8_32_29_inst0__config_addr[7:0] = config_config_addr[7:0];

  assign ConfigRegister_1_8_32_29_inst0__config_data[31:0] = config_config_data[31:0];

  assign ConfigRegister_1_8_32_29_inst0__config_en = config_write[0];

  assign ConfigRegister_1_8_32_29_inst0__reset = reset;

  assign MuxWrapper_2_16_inst5__S[0:0] = ConfigRegister_1_8_32_31_inst0__O[0:0];

  assign ZextWrapper_1_32_inst15__I[0:0] = ConfigRegister_1_8_32_31_inst0__O[0:0];

  assign ConfigRegister_1_8_32_31_inst0__clk = clk;

  assign ConfigRegister_1_8_32_31_inst0__config_addr[7:0] = config_config_addr[7:0];

  assign ConfigRegister_1_8_32_31_inst0__config_data[31:0] = config_config_data[31:0];

  assign ConfigRegister_1_8_32_31_inst0__config_en = config_write[0];

  assign ConfigRegister_1_8_32_31_inst0__reset = reset;

  assign MuxWrapper_2_16_inst6__S[0:0] = ConfigRegister_1_8_32_33_inst0__O[0:0];

  assign ZextWrapper_1_32_inst16__I[0:0] = ConfigRegister_1_8_32_33_inst0__O[0:0];

  assign ConfigRegister_1_8_32_33_inst0__clk = clk;

  assign ConfigRegister_1_8_32_33_inst0__config_addr[7:0] = config_config_addr[7:0];

  assign ConfigRegister_1_8_32_33_inst0__config_data[31:0] = config_config_data[31:0];

  assign ConfigRegister_1_8_32_33_inst0__config_en = config_write[0];

  assign ConfigRegister_1_8_32_33_inst0__reset = reset;

  assign MuxWrapper_2_16_inst7__S[0:0] = ConfigRegister_1_8_32_35_inst0__O[0:0];

  assign ZextWrapper_1_32_inst17__I[0:0] = ConfigRegister_1_8_32_35_inst0__O[0:0];

  assign ConfigRegister_1_8_32_35_inst0__clk = clk;

  assign ConfigRegister_1_8_32_35_inst0__config_addr[7:0] = config_config_addr[7:0];

  assign ConfigRegister_1_8_32_35_inst0__config_data[31:0] = config_config_data[31:0];

  assign ConfigRegister_1_8_32_35_inst0__config_en = config_write[0];

  assign ConfigRegister_1_8_32_35_inst0__reset = reset;

  assign MuxWrapper_2_16_inst8__S[0:0] = ConfigRegister_1_8_32_37_inst0__O[0:0];

  assign ZextWrapper_1_32_inst18__I[0:0] = ConfigRegister_1_8_32_37_inst0__O[0:0];

  assign ConfigRegister_1_8_32_37_inst0__clk = clk;

  assign ConfigRegister_1_8_32_37_inst0__config_addr[7:0] = config_config_addr[7:0];

  assign ConfigRegister_1_8_32_37_inst0__config_data[31:0] = config_config_data[31:0];

  assign ConfigRegister_1_8_32_37_inst0__config_en = config_write[0];

  assign ConfigRegister_1_8_32_37_inst0__reset = reset;

  assign MuxWrapper_2_16_inst9__S[0:0] = ConfigRegister_1_8_32_39_inst0__O[0:0];

  assign ZextWrapper_1_32_inst19__I[0:0] = ConfigRegister_1_8_32_39_inst0__O[0:0];

  assign ConfigRegister_1_8_32_39_inst0__clk = clk;

  assign ConfigRegister_1_8_32_39_inst0__config_addr[7:0] = config_config_addr[7:0];

  assign ConfigRegister_1_8_32_39_inst0__config_data[31:0] = config_config_data[31:0];

  assign ConfigRegister_1_8_32_39_inst0__config_en = config_write[0];

  assign ConfigRegister_1_8_32_39_inst0__reset = reset;

  assign MuxWrapper_2_1_inst1__S[0:0] = ConfigRegister_1_8_32_3_inst0__O[0:0];

  assign ZextWrapper_1_32_inst1__I[0:0] = ConfigRegister_1_8_32_3_inst0__O[0:0];

  assign ConfigRegister_1_8_32_3_inst0__clk = clk;

  assign ConfigRegister_1_8_32_3_inst0__config_addr[7:0] = config_config_addr[7:0];

  assign ConfigRegister_1_8_32_3_inst0__config_data[31:0] = config_config_data[31:0];

  assign ConfigRegister_1_8_32_3_inst0__config_en = config_write[0];

  assign ConfigRegister_1_8_32_3_inst0__reset = reset;

  assign MuxWrapper_2_1_inst10__S[0:0] = ConfigRegister_1_8_32_41_inst0__O[0:0];

  assign ZextWrapper_1_32_inst20__I[0:0] = ConfigRegister_1_8_32_41_inst0__O[0:0];

  assign ConfigRegister_1_8_32_41_inst0__clk = clk;

  assign ConfigRegister_1_8_32_41_inst0__config_addr[7:0] = config_config_addr[7:0];

  assign ConfigRegister_1_8_32_41_inst0__config_data[31:0] = config_config_data[31:0];

  assign ConfigRegister_1_8_32_41_inst0__config_en = config_write[0];

  assign ConfigRegister_1_8_32_41_inst0__reset = reset;

  assign MuxWrapper_2_1_inst11__S[0:0] = ConfigRegister_1_8_32_43_inst0__O[0:0];

  assign ZextWrapper_1_32_inst21__I[0:0] = ConfigRegister_1_8_32_43_inst0__O[0:0];

  assign ConfigRegister_1_8_32_43_inst0__clk = clk;

  assign ConfigRegister_1_8_32_43_inst0__config_addr[7:0] = config_config_addr[7:0];

  assign ConfigRegister_1_8_32_43_inst0__config_data[31:0] = config_config_data[31:0];

  assign ConfigRegister_1_8_32_43_inst0__config_en = config_write[0];

  assign ConfigRegister_1_8_32_43_inst0__reset = reset;

  assign MuxWrapper_2_1_inst12__S[0:0] = ConfigRegister_1_8_32_45_inst0__O[0:0];

  assign ZextWrapper_1_32_inst22__I[0:0] = ConfigRegister_1_8_32_45_inst0__O[0:0];

  assign ConfigRegister_1_8_32_45_inst0__clk = clk;

  assign ConfigRegister_1_8_32_45_inst0__config_addr[7:0] = config_config_addr[7:0];

  assign ConfigRegister_1_8_32_45_inst0__config_data[31:0] = config_config_data[31:0];

  assign ConfigRegister_1_8_32_45_inst0__config_en = config_write[0];

  assign ConfigRegister_1_8_32_45_inst0__reset = reset;

  assign MuxWrapper_2_1_inst13__S[0:0] = ConfigRegister_1_8_32_47_inst0__O[0:0];

  assign ZextWrapper_1_32_inst23__I[0:0] = ConfigRegister_1_8_32_47_inst0__O[0:0];

  assign ConfigRegister_1_8_32_47_inst0__clk = clk;

  assign ConfigRegister_1_8_32_47_inst0__config_addr[7:0] = config_config_addr[7:0];

  assign ConfigRegister_1_8_32_47_inst0__config_data[31:0] = config_config_data[31:0];

  assign ConfigRegister_1_8_32_47_inst0__config_en = config_write[0];

  assign ConfigRegister_1_8_32_47_inst0__reset = reset;

  assign MuxWrapper_2_1_inst14__S[0:0] = ConfigRegister_1_8_32_49_inst0__O[0:0];

  assign ZextWrapper_1_32_inst24__I[0:0] = ConfigRegister_1_8_32_49_inst0__O[0:0];

  assign ConfigRegister_1_8_32_49_inst0__clk = clk;

  assign ConfigRegister_1_8_32_49_inst0__config_addr[7:0] = config_config_addr[7:0];

  assign ConfigRegister_1_8_32_49_inst0__config_data[31:0] = config_config_data[31:0];

  assign ConfigRegister_1_8_32_49_inst0__config_en = config_write[0];

  assign ConfigRegister_1_8_32_49_inst0__reset = reset;

  assign MuxWrapper_2_16_inst10__S[0:0] = ConfigRegister_1_8_32_51_inst0__O[0:0];

  assign ZextWrapper_1_32_inst25__I[0:0] = ConfigRegister_1_8_32_51_inst0__O[0:0];

  assign ConfigRegister_1_8_32_51_inst0__clk = clk;

  assign ConfigRegister_1_8_32_51_inst0__config_addr[7:0] = config_config_addr[7:0];

  assign ConfigRegister_1_8_32_51_inst0__config_data[31:0] = config_config_data[31:0];

  assign ConfigRegister_1_8_32_51_inst0__config_en = config_write[0];

  assign ConfigRegister_1_8_32_51_inst0__reset = reset;

  assign MuxWrapper_2_16_inst11__S[0:0] = ConfigRegister_1_8_32_53_inst0__O[0:0];

  assign ZextWrapper_1_32_inst26__I[0:0] = ConfigRegister_1_8_32_53_inst0__O[0:0];

  assign ConfigRegister_1_8_32_53_inst0__clk = clk;

  assign ConfigRegister_1_8_32_53_inst0__config_addr[7:0] = config_config_addr[7:0];

  assign ConfigRegister_1_8_32_53_inst0__config_data[31:0] = config_config_data[31:0];

  assign ConfigRegister_1_8_32_53_inst0__config_en = config_write[0];

  assign ConfigRegister_1_8_32_53_inst0__reset = reset;

  assign MuxWrapper_2_16_inst12__S[0:0] = ConfigRegister_1_8_32_55_inst0__O[0:0];

  assign ZextWrapper_1_32_inst27__I[0:0] = ConfigRegister_1_8_32_55_inst0__O[0:0];

  assign ConfigRegister_1_8_32_55_inst0__clk = clk;

  assign ConfigRegister_1_8_32_55_inst0__config_addr[7:0] = config_config_addr[7:0];

  assign ConfigRegister_1_8_32_55_inst0__config_data[31:0] = config_config_data[31:0];

  assign ConfigRegister_1_8_32_55_inst0__config_en = config_write[0];

  assign ConfigRegister_1_8_32_55_inst0__reset = reset;

  assign MuxWrapper_2_16_inst13__S[0:0] = ConfigRegister_1_8_32_57_inst0__O[0:0];

  assign ZextWrapper_1_32_inst28__I[0:0] = ConfigRegister_1_8_32_57_inst0__O[0:0];

  assign ConfigRegister_1_8_32_57_inst0__clk = clk;

  assign ConfigRegister_1_8_32_57_inst0__config_addr[7:0] = config_config_addr[7:0];

  assign ConfigRegister_1_8_32_57_inst0__config_data[31:0] = config_config_data[31:0];

  assign ConfigRegister_1_8_32_57_inst0__config_en = config_write[0];

  assign ConfigRegister_1_8_32_57_inst0__reset = reset;

  assign MuxWrapper_2_16_inst14__S[0:0] = ConfigRegister_1_8_32_59_inst0__O[0:0];

  assign ZextWrapper_1_32_inst29__I[0:0] = ConfigRegister_1_8_32_59_inst0__O[0:0];

  assign ConfigRegister_1_8_32_59_inst0__clk = clk;

  assign ConfigRegister_1_8_32_59_inst0__config_addr[7:0] = config_config_addr[7:0];

  assign ConfigRegister_1_8_32_59_inst0__config_data[31:0] = config_config_data[31:0];

  assign ConfigRegister_1_8_32_59_inst0__config_en = config_write[0];

  assign ConfigRegister_1_8_32_59_inst0__reset = reset;

  assign MuxWrapper_2_1_inst2__S[0:0] = ConfigRegister_1_8_32_5_inst0__O[0:0];

  assign ZextWrapper_1_32_inst2__I[0:0] = ConfigRegister_1_8_32_5_inst0__O[0:0];

  assign ConfigRegister_1_8_32_5_inst0__clk = clk;

  assign ConfigRegister_1_8_32_5_inst0__config_addr[7:0] = config_config_addr[7:0];

  assign ConfigRegister_1_8_32_5_inst0__config_data[31:0] = config_config_data[31:0];

  assign ConfigRegister_1_8_32_5_inst0__config_en = config_write[0];

  assign ConfigRegister_1_8_32_5_inst0__reset = reset;

  assign MuxWrapper_2_1_inst15__S[0:0] = ConfigRegister_1_8_32_61_inst0__O[0:0];

  assign ZextWrapper_1_32_inst30__I[0:0] = ConfigRegister_1_8_32_61_inst0__O[0:0];

  assign ConfigRegister_1_8_32_61_inst0__clk = clk;

  assign ConfigRegister_1_8_32_61_inst0__config_addr[7:0] = config_config_addr[7:0];

  assign ConfigRegister_1_8_32_61_inst0__config_data[31:0] = config_config_data[31:0];

  assign ConfigRegister_1_8_32_61_inst0__config_en = config_write[0];

  assign ConfigRegister_1_8_32_61_inst0__reset = reset;

  assign MuxWrapper_2_1_inst16__S[0:0] = ConfigRegister_1_8_32_63_inst0__O[0:0];

  assign ZextWrapper_1_32_inst31__I[0:0] = ConfigRegister_1_8_32_63_inst0__O[0:0];

  assign ConfigRegister_1_8_32_63_inst0__clk = clk;

  assign ConfigRegister_1_8_32_63_inst0__config_addr[7:0] = config_config_addr[7:0];

  assign ConfigRegister_1_8_32_63_inst0__config_data[31:0] = config_config_data[31:0];

  assign ConfigRegister_1_8_32_63_inst0__config_en = config_write[0];

  assign ConfigRegister_1_8_32_63_inst0__reset = reset;

  assign MuxWrapper_2_1_inst17__S[0:0] = ConfigRegister_1_8_32_65_inst0__O[0:0];

  assign ZextWrapper_1_32_inst32__I[0:0] = ConfigRegister_1_8_32_65_inst0__O[0:0];

  assign ConfigRegister_1_8_32_65_inst0__clk = clk;

  assign ConfigRegister_1_8_32_65_inst0__config_addr[7:0] = config_config_addr[7:0];

  assign ConfigRegister_1_8_32_65_inst0__config_data[31:0] = config_config_data[31:0];

  assign ConfigRegister_1_8_32_65_inst0__config_en = config_write[0];

  assign ConfigRegister_1_8_32_65_inst0__reset = reset;

  assign MuxWrapper_2_1_inst18__S[0:0] = ConfigRegister_1_8_32_67_inst0__O[0:0];

  assign ZextWrapper_1_32_inst33__I[0:0] = ConfigRegister_1_8_32_67_inst0__O[0:0];

  assign ConfigRegister_1_8_32_67_inst0__clk = clk;

  assign ConfigRegister_1_8_32_67_inst0__config_addr[7:0] = config_config_addr[7:0];

  assign ConfigRegister_1_8_32_67_inst0__config_data[31:0] = config_config_data[31:0];

  assign ConfigRegister_1_8_32_67_inst0__config_en = config_write[0];

  assign ConfigRegister_1_8_32_67_inst0__reset = reset;

  assign MuxWrapper_2_1_inst19__S[0:0] = ConfigRegister_1_8_32_69_inst0__O[0:0];

  assign ZextWrapper_1_32_inst34__I[0:0] = ConfigRegister_1_8_32_69_inst0__O[0:0];

  assign ConfigRegister_1_8_32_69_inst0__clk = clk;

  assign ConfigRegister_1_8_32_69_inst0__config_addr[7:0] = config_config_addr[7:0];

  assign ConfigRegister_1_8_32_69_inst0__config_data[31:0] = config_config_data[31:0];

  assign ConfigRegister_1_8_32_69_inst0__config_en = config_write[0];

  assign ConfigRegister_1_8_32_69_inst0__reset = reset;

  assign MuxWrapper_2_16_inst15__S[0:0] = ConfigRegister_1_8_32_71_inst0__O[0:0];

  assign ZextWrapper_1_32_inst35__I[0:0] = ConfigRegister_1_8_32_71_inst0__O[0:0];

  assign ConfigRegister_1_8_32_71_inst0__clk = clk;

  assign ConfigRegister_1_8_32_71_inst0__config_addr[7:0] = config_config_addr[7:0];

  assign ConfigRegister_1_8_32_71_inst0__config_data[31:0] = config_config_data[31:0];

  assign ConfigRegister_1_8_32_71_inst0__config_en = config_write[0];

  assign ConfigRegister_1_8_32_71_inst0__reset = reset;

  assign MuxWrapper_2_16_inst16__S[0:0] = ConfigRegister_1_8_32_73_inst0__O[0:0];

  assign ZextWrapper_1_32_inst36__I[0:0] = ConfigRegister_1_8_32_73_inst0__O[0:0];

  assign ConfigRegister_1_8_32_73_inst0__clk = clk;

  assign ConfigRegister_1_8_32_73_inst0__config_addr[7:0] = config_config_addr[7:0];

  assign ConfigRegister_1_8_32_73_inst0__config_data[31:0] = config_config_data[31:0];

  assign ConfigRegister_1_8_32_73_inst0__config_en = config_write[0];

  assign ConfigRegister_1_8_32_73_inst0__reset = reset;

  assign MuxWrapper_2_16_inst17__S[0:0] = ConfigRegister_1_8_32_75_inst0__O[0:0];

  assign ZextWrapper_1_32_inst37__I[0:0] = ConfigRegister_1_8_32_75_inst0__O[0:0];

  assign ConfigRegister_1_8_32_75_inst0__clk = clk;

  assign ConfigRegister_1_8_32_75_inst0__config_addr[7:0] = config_config_addr[7:0];

  assign ConfigRegister_1_8_32_75_inst0__config_data[31:0] = config_config_data[31:0];

  assign ConfigRegister_1_8_32_75_inst0__config_en = config_write[0];

  assign ConfigRegister_1_8_32_75_inst0__reset = reset;

  assign MuxWrapper_2_16_inst18__S[0:0] = ConfigRegister_1_8_32_77_inst0__O[0:0];

  assign ZextWrapper_1_32_inst38__I[0:0] = ConfigRegister_1_8_32_77_inst0__O[0:0];

  assign ConfigRegister_1_8_32_77_inst0__clk = clk;

  assign ConfigRegister_1_8_32_77_inst0__config_addr[7:0] = config_config_addr[7:0];

  assign ConfigRegister_1_8_32_77_inst0__config_data[31:0] = config_config_data[31:0];

  assign ConfigRegister_1_8_32_77_inst0__config_en = config_write[0];

  assign ConfigRegister_1_8_32_77_inst0__reset = reset;

  assign MuxWrapper_2_16_inst19__S[0:0] = ConfigRegister_1_8_32_79_inst0__O[0:0];

  assign ZextWrapper_1_32_inst39__I[0:0] = ConfigRegister_1_8_32_79_inst0__O[0:0];

  assign ConfigRegister_1_8_32_79_inst0__clk = clk;

  assign ConfigRegister_1_8_32_79_inst0__config_addr[7:0] = config_config_addr[7:0];

  assign ConfigRegister_1_8_32_79_inst0__config_data[31:0] = config_config_data[31:0];

  assign ConfigRegister_1_8_32_79_inst0__config_en = config_write[0];

  assign ConfigRegister_1_8_32_79_inst0__reset = reset;

  assign MuxWrapper_2_1_inst3__S[0:0] = ConfigRegister_1_8_32_7_inst0__O[0:0];

  assign ZextWrapper_1_32_inst3__I[0:0] = ConfigRegister_1_8_32_7_inst0__O[0:0];

  assign ConfigRegister_1_8_32_7_inst0__clk = clk;

  assign ConfigRegister_1_8_32_7_inst0__config_addr[7:0] = config_config_addr[7:0];

  assign ConfigRegister_1_8_32_7_inst0__config_data[31:0] = config_config_data[31:0];

  assign ConfigRegister_1_8_32_7_inst0__config_en = config_write[0];

  assign ConfigRegister_1_8_32_7_inst0__reset = reset;

  assign MuxWrapper_2_1_inst4__S[0:0] = ConfigRegister_1_8_32_9_inst0__O[0:0];

  assign ZextWrapper_1_32_inst4__I[0:0] = ConfigRegister_1_8_32_9_inst0__O[0:0];

  assign ConfigRegister_1_8_32_9_inst0__clk = clk;

  assign ConfigRegister_1_8_32_9_inst0__config_addr[7:0] = config_config_addr[7:0];

  assign ConfigRegister_1_8_32_9_inst0__config_data[31:0] = config_config_data[31:0];

  assign ConfigRegister_1_8_32_9_inst0__config_en = config_write[0];

  assign ConfigRegister_1_8_32_9_inst0__reset = reset;

  assign MuxWrapper_4_1_inst0__S[1:0] = ConfigRegister_2_8_32_0_inst0__O[1:0];

  assign ZextWrapper_2_32_inst0__I[1:0] = ConfigRegister_2_8_32_0_inst0__O[1:0];

  assign ConfigRegister_2_8_32_0_inst0__clk = clk;

  assign ConfigRegister_2_8_32_0_inst0__config_addr[7:0] = config_config_addr[7:0];

  assign ConfigRegister_2_8_32_0_inst0__config_data[31:0] = config_config_data[31:0];

  assign ConfigRegister_2_8_32_0_inst0__config_en = config_write[0];

  assign ConfigRegister_2_8_32_0_inst0__reset = reset;

  assign MuxWrapper_4_16_inst0__S[1:0] = ConfigRegister_2_8_32_10_inst0__O[1:0];

  assign ZextWrapper_2_32_inst5__I[1:0] = ConfigRegister_2_8_32_10_inst0__O[1:0];

  assign ConfigRegister_2_8_32_10_inst0__clk = clk;

  assign ConfigRegister_2_8_32_10_inst0__config_addr[7:0] = config_config_addr[7:0];

  assign ConfigRegister_2_8_32_10_inst0__config_data[31:0] = config_config_data[31:0];

  assign ConfigRegister_2_8_32_10_inst0__config_en = config_write[0];

  assign ConfigRegister_2_8_32_10_inst0__reset = reset;

  assign MuxWrapper_4_16_inst1__S[1:0] = ConfigRegister_2_8_32_12_inst0__O[1:0];

  assign ZextWrapper_2_32_inst6__I[1:0] = ConfigRegister_2_8_32_12_inst0__O[1:0];

  assign ConfigRegister_2_8_32_12_inst0__clk = clk;

  assign ConfigRegister_2_8_32_12_inst0__config_addr[7:0] = config_config_addr[7:0];

  assign ConfigRegister_2_8_32_12_inst0__config_data[31:0] = config_config_data[31:0];

  assign ConfigRegister_2_8_32_12_inst0__config_en = config_write[0];

  assign ConfigRegister_2_8_32_12_inst0__reset = reset;

  assign MuxWrapper_4_16_inst2__S[1:0] = ConfigRegister_2_8_32_14_inst0__O[1:0];

  assign ZextWrapper_2_32_inst7__I[1:0] = ConfigRegister_2_8_32_14_inst0__O[1:0];

  assign ConfigRegister_2_8_32_14_inst0__clk = clk;

  assign ConfigRegister_2_8_32_14_inst0__config_addr[7:0] = config_config_addr[7:0];

  assign ConfigRegister_2_8_32_14_inst0__config_data[31:0] = config_config_data[31:0];

  assign ConfigRegister_2_8_32_14_inst0__config_en = config_write[0];

  assign ConfigRegister_2_8_32_14_inst0__reset = reset;

  assign MuxWrapper_4_16_inst3__S[1:0] = ConfigRegister_2_8_32_16_inst0__O[1:0];

  assign ZextWrapper_2_32_inst8__I[1:0] = ConfigRegister_2_8_32_16_inst0__O[1:0];

  assign ConfigRegister_2_8_32_16_inst0__clk = clk;

  assign ConfigRegister_2_8_32_16_inst0__config_addr[7:0] = config_config_addr[7:0];

  assign ConfigRegister_2_8_32_16_inst0__config_data[31:0] = config_config_data[31:0];

  assign ConfigRegister_2_8_32_16_inst0__config_en = config_write[0];

  assign ConfigRegister_2_8_32_16_inst0__reset = reset;

  assign MuxWrapper_4_16_inst4__S[1:0] = ConfigRegister_2_8_32_18_inst0__O[1:0];

  assign ZextWrapper_2_32_inst9__I[1:0] = ConfigRegister_2_8_32_18_inst0__O[1:0];

  assign ConfigRegister_2_8_32_18_inst0__clk = clk;

  assign ConfigRegister_2_8_32_18_inst0__config_addr[7:0] = config_config_addr[7:0];

  assign ConfigRegister_2_8_32_18_inst0__config_data[31:0] = config_config_data[31:0];

  assign ConfigRegister_2_8_32_18_inst0__config_en = config_write[0];

  assign ConfigRegister_2_8_32_18_inst0__reset = reset;

  assign MuxWrapper_4_1_inst5__S[1:0] = ConfigRegister_2_8_32_20_inst0__O[1:0];

  assign ZextWrapper_2_32_inst10__I[1:0] = ConfigRegister_2_8_32_20_inst0__O[1:0];

  assign ConfigRegister_2_8_32_20_inst0__clk = clk;

  assign ConfigRegister_2_8_32_20_inst0__config_addr[7:0] = config_config_addr[7:0];

  assign ConfigRegister_2_8_32_20_inst0__config_data[31:0] = config_config_data[31:0];

  assign ConfigRegister_2_8_32_20_inst0__config_en = config_write[0];

  assign ConfigRegister_2_8_32_20_inst0__reset = reset;

  assign MuxWrapper_4_1_inst6__S[1:0] = ConfigRegister_2_8_32_22_inst0__O[1:0];

  assign ZextWrapper_2_32_inst11__I[1:0] = ConfigRegister_2_8_32_22_inst0__O[1:0];

  assign ConfigRegister_2_8_32_22_inst0__clk = clk;

  assign ConfigRegister_2_8_32_22_inst0__config_addr[7:0] = config_config_addr[7:0];

  assign ConfigRegister_2_8_32_22_inst0__config_data[31:0] = config_config_data[31:0];

  assign ConfigRegister_2_8_32_22_inst0__config_en = config_write[0];

  assign ConfigRegister_2_8_32_22_inst0__reset = reset;

  assign MuxWrapper_4_1_inst7__S[1:0] = ConfigRegister_2_8_32_24_inst0__O[1:0];

  assign ZextWrapper_2_32_inst12__I[1:0] = ConfigRegister_2_8_32_24_inst0__O[1:0];

  assign ConfigRegister_2_8_32_24_inst0__clk = clk;

  assign ConfigRegister_2_8_32_24_inst0__config_addr[7:0] = config_config_addr[7:0];

  assign ConfigRegister_2_8_32_24_inst0__config_data[31:0] = config_config_data[31:0];

  assign ConfigRegister_2_8_32_24_inst0__config_en = config_write[0];

  assign ConfigRegister_2_8_32_24_inst0__reset = reset;

  assign MuxWrapper_4_1_inst8__S[1:0] = ConfigRegister_2_8_32_26_inst0__O[1:0];

  assign ZextWrapper_2_32_inst13__I[1:0] = ConfigRegister_2_8_32_26_inst0__O[1:0];

  assign ConfigRegister_2_8_32_26_inst0__clk = clk;

  assign ConfigRegister_2_8_32_26_inst0__config_addr[7:0] = config_config_addr[7:0];

  assign ConfigRegister_2_8_32_26_inst0__config_data[31:0] = config_config_data[31:0];

  assign ConfigRegister_2_8_32_26_inst0__config_en = config_write[0];

  assign ConfigRegister_2_8_32_26_inst0__reset = reset;

  assign MuxWrapper_4_1_inst9__S[1:0] = ConfigRegister_2_8_32_28_inst0__O[1:0];

  assign ZextWrapper_2_32_inst14__I[1:0] = ConfigRegister_2_8_32_28_inst0__O[1:0];

  assign ConfigRegister_2_8_32_28_inst0__clk = clk;

  assign ConfigRegister_2_8_32_28_inst0__config_addr[7:0] = config_config_addr[7:0];

  assign ConfigRegister_2_8_32_28_inst0__config_data[31:0] = config_config_data[31:0];

  assign ConfigRegister_2_8_32_28_inst0__config_en = config_write[0];

  assign ConfigRegister_2_8_32_28_inst0__reset = reset;

  assign MuxWrapper_4_1_inst1__S[1:0] = ConfigRegister_2_8_32_2_inst0__O[1:0];

  assign ZextWrapper_2_32_inst1__I[1:0] = ConfigRegister_2_8_32_2_inst0__O[1:0];

  assign ConfigRegister_2_8_32_2_inst0__clk = clk;

  assign ConfigRegister_2_8_32_2_inst0__config_addr[7:0] = config_config_addr[7:0];

  assign ConfigRegister_2_8_32_2_inst0__config_data[31:0] = config_config_data[31:0];

  assign ConfigRegister_2_8_32_2_inst0__config_en = config_write[0];

  assign ConfigRegister_2_8_32_2_inst0__reset = reset;

  assign MuxWrapper_4_16_inst5__S[1:0] = ConfigRegister_2_8_32_30_inst0__O[1:0];

  assign ZextWrapper_2_32_inst15__I[1:0] = ConfigRegister_2_8_32_30_inst0__O[1:0];

  assign ConfigRegister_2_8_32_30_inst0__clk = clk;

  assign ConfigRegister_2_8_32_30_inst0__config_addr[7:0] = config_config_addr[7:0];

  assign ConfigRegister_2_8_32_30_inst0__config_data[31:0] = config_config_data[31:0];

  assign ConfigRegister_2_8_32_30_inst0__config_en = config_write[0];

  assign ConfigRegister_2_8_32_30_inst0__reset = reset;

  assign MuxWrapper_4_16_inst6__S[1:0] = ConfigRegister_2_8_32_32_inst0__O[1:0];

  assign ZextWrapper_2_32_inst16__I[1:0] = ConfigRegister_2_8_32_32_inst0__O[1:0];

  assign ConfigRegister_2_8_32_32_inst0__clk = clk;

  assign ConfigRegister_2_8_32_32_inst0__config_addr[7:0] = config_config_addr[7:0];

  assign ConfigRegister_2_8_32_32_inst0__config_data[31:0] = config_config_data[31:0];

  assign ConfigRegister_2_8_32_32_inst0__config_en = config_write[0];

  assign ConfigRegister_2_8_32_32_inst0__reset = reset;

  assign MuxWrapper_4_16_inst7__S[1:0] = ConfigRegister_2_8_32_34_inst0__O[1:0];

  assign ZextWrapper_2_32_inst17__I[1:0] = ConfigRegister_2_8_32_34_inst0__O[1:0];

  assign ConfigRegister_2_8_32_34_inst0__clk = clk;

  assign ConfigRegister_2_8_32_34_inst0__config_addr[7:0] = config_config_addr[7:0];

  assign ConfigRegister_2_8_32_34_inst0__config_data[31:0] = config_config_data[31:0];

  assign ConfigRegister_2_8_32_34_inst0__config_en = config_write[0];

  assign ConfigRegister_2_8_32_34_inst0__reset = reset;

  assign MuxWrapper_4_16_inst8__S[1:0] = ConfigRegister_2_8_32_36_inst0__O[1:0];

  assign ZextWrapper_2_32_inst18__I[1:0] = ConfigRegister_2_8_32_36_inst0__O[1:0];

  assign ConfigRegister_2_8_32_36_inst0__clk = clk;

  assign ConfigRegister_2_8_32_36_inst0__config_addr[7:0] = config_config_addr[7:0];

  assign ConfigRegister_2_8_32_36_inst0__config_data[31:0] = config_config_data[31:0];

  assign ConfigRegister_2_8_32_36_inst0__config_en = config_write[0];

  assign ConfigRegister_2_8_32_36_inst0__reset = reset;

  assign MuxWrapper_4_16_inst9__S[1:0] = ConfigRegister_2_8_32_38_inst0__O[1:0];

  assign ZextWrapper_2_32_inst19__I[1:0] = ConfigRegister_2_8_32_38_inst0__O[1:0];

  assign ConfigRegister_2_8_32_38_inst0__clk = clk;

  assign ConfigRegister_2_8_32_38_inst0__config_addr[7:0] = config_config_addr[7:0];

  assign ConfigRegister_2_8_32_38_inst0__config_data[31:0] = config_config_data[31:0];

  assign ConfigRegister_2_8_32_38_inst0__config_en = config_write[0];

  assign ConfigRegister_2_8_32_38_inst0__reset = reset;

  assign MuxWrapper_4_1_inst10__S[1:0] = ConfigRegister_2_8_32_40_inst0__O[1:0];

  assign ZextWrapper_2_32_inst20__I[1:0] = ConfigRegister_2_8_32_40_inst0__O[1:0];

  assign ConfigRegister_2_8_32_40_inst0__clk = clk;

  assign ConfigRegister_2_8_32_40_inst0__config_addr[7:0] = config_config_addr[7:0];

  assign ConfigRegister_2_8_32_40_inst0__config_data[31:0] = config_config_data[31:0];

  assign ConfigRegister_2_8_32_40_inst0__config_en = config_write[0];

  assign ConfigRegister_2_8_32_40_inst0__reset = reset;

  assign MuxWrapper_4_1_inst11__S[1:0] = ConfigRegister_2_8_32_42_inst0__O[1:0];

  assign ZextWrapper_2_32_inst21__I[1:0] = ConfigRegister_2_8_32_42_inst0__O[1:0];

  assign ConfigRegister_2_8_32_42_inst0__clk = clk;

  assign ConfigRegister_2_8_32_42_inst0__config_addr[7:0] = config_config_addr[7:0];

  assign ConfigRegister_2_8_32_42_inst0__config_data[31:0] = config_config_data[31:0];

  assign ConfigRegister_2_8_32_42_inst0__config_en = config_write[0];

  assign ConfigRegister_2_8_32_42_inst0__reset = reset;

  assign MuxWrapper_4_1_inst12__S[1:0] = ConfigRegister_2_8_32_44_inst0__O[1:0];

  assign ZextWrapper_2_32_inst22__I[1:0] = ConfigRegister_2_8_32_44_inst0__O[1:0];

  assign ConfigRegister_2_8_32_44_inst0__clk = clk;

  assign ConfigRegister_2_8_32_44_inst0__config_addr[7:0] = config_config_addr[7:0];

  assign ConfigRegister_2_8_32_44_inst0__config_data[31:0] = config_config_data[31:0];

  assign ConfigRegister_2_8_32_44_inst0__config_en = config_write[0];

  assign ConfigRegister_2_8_32_44_inst0__reset = reset;

  assign MuxWrapper_4_1_inst13__S[1:0] = ConfigRegister_2_8_32_46_inst0__O[1:0];

  assign ZextWrapper_2_32_inst23__I[1:0] = ConfigRegister_2_8_32_46_inst0__O[1:0];

  assign ConfigRegister_2_8_32_46_inst0__clk = clk;

  assign ConfigRegister_2_8_32_46_inst0__config_addr[7:0] = config_config_addr[7:0];

  assign ConfigRegister_2_8_32_46_inst0__config_data[31:0] = config_config_data[31:0];

  assign ConfigRegister_2_8_32_46_inst0__config_en = config_write[0];

  assign ConfigRegister_2_8_32_46_inst0__reset = reset;

  assign MuxWrapper_4_1_inst14__S[1:0] = ConfigRegister_2_8_32_48_inst0__O[1:0];

  assign ZextWrapper_2_32_inst24__I[1:0] = ConfigRegister_2_8_32_48_inst0__O[1:0];

  assign ConfigRegister_2_8_32_48_inst0__clk = clk;

  assign ConfigRegister_2_8_32_48_inst0__config_addr[7:0] = config_config_addr[7:0];

  assign ConfigRegister_2_8_32_48_inst0__config_data[31:0] = config_config_data[31:0];

  assign ConfigRegister_2_8_32_48_inst0__config_en = config_write[0];

  assign ConfigRegister_2_8_32_48_inst0__reset = reset;

  assign MuxWrapper_4_1_inst2__S[1:0] = ConfigRegister_2_8_32_4_inst0__O[1:0];

  assign ZextWrapper_2_32_inst2__I[1:0] = ConfigRegister_2_8_32_4_inst0__O[1:0];

  assign ConfigRegister_2_8_32_4_inst0__clk = clk;

  assign ConfigRegister_2_8_32_4_inst0__config_addr[7:0] = config_config_addr[7:0];

  assign ConfigRegister_2_8_32_4_inst0__config_data[31:0] = config_config_data[31:0];

  assign ConfigRegister_2_8_32_4_inst0__config_en = config_write[0];

  assign ConfigRegister_2_8_32_4_inst0__reset = reset;

  assign MuxWrapper_4_16_inst10__S[1:0] = ConfigRegister_2_8_32_50_inst0__O[1:0];

  assign ZextWrapper_2_32_inst25__I[1:0] = ConfigRegister_2_8_32_50_inst0__O[1:0];

  assign ConfigRegister_2_8_32_50_inst0__clk = clk;

  assign ConfigRegister_2_8_32_50_inst0__config_addr[7:0] = config_config_addr[7:0];

  assign ConfigRegister_2_8_32_50_inst0__config_data[31:0] = config_config_data[31:0];

  assign ConfigRegister_2_8_32_50_inst0__config_en = config_write[0];

  assign ConfigRegister_2_8_32_50_inst0__reset = reset;

  assign MuxWrapper_4_16_inst11__S[1:0] = ConfigRegister_2_8_32_52_inst0__O[1:0];

  assign ZextWrapper_2_32_inst26__I[1:0] = ConfigRegister_2_8_32_52_inst0__O[1:0];

  assign ConfigRegister_2_8_32_52_inst0__clk = clk;

  assign ConfigRegister_2_8_32_52_inst0__config_addr[7:0] = config_config_addr[7:0];

  assign ConfigRegister_2_8_32_52_inst0__config_data[31:0] = config_config_data[31:0];

  assign ConfigRegister_2_8_32_52_inst0__config_en = config_write[0];

  assign ConfigRegister_2_8_32_52_inst0__reset = reset;

  assign MuxWrapper_4_16_inst12__S[1:0] = ConfigRegister_2_8_32_54_inst0__O[1:0];

  assign ZextWrapper_2_32_inst27__I[1:0] = ConfigRegister_2_8_32_54_inst0__O[1:0];

  assign ConfigRegister_2_8_32_54_inst0__clk = clk;

  assign ConfigRegister_2_8_32_54_inst0__config_addr[7:0] = config_config_addr[7:0];

  assign ConfigRegister_2_8_32_54_inst0__config_data[31:0] = config_config_data[31:0];

  assign ConfigRegister_2_8_32_54_inst0__config_en = config_write[0];

  assign ConfigRegister_2_8_32_54_inst0__reset = reset;

  assign MuxWrapper_4_16_inst13__S[1:0] = ConfigRegister_2_8_32_56_inst0__O[1:0];

  assign ZextWrapper_2_32_inst28__I[1:0] = ConfigRegister_2_8_32_56_inst0__O[1:0];

  assign ConfigRegister_2_8_32_56_inst0__clk = clk;

  assign ConfigRegister_2_8_32_56_inst0__config_addr[7:0] = config_config_addr[7:0];

  assign ConfigRegister_2_8_32_56_inst0__config_data[31:0] = config_config_data[31:0];

  assign ConfigRegister_2_8_32_56_inst0__config_en = config_write[0];

  assign ConfigRegister_2_8_32_56_inst0__reset = reset;

  assign MuxWrapper_4_16_inst14__S[1:0] = ConfigRegister_2_8_32_58_inst0__O[1:0];

  assign ZextWrapper_2_32_inst29__I[1:0] = ConfigRegister_2_8_32_58_inst0__O[1:0];

  assign ConfigRegister_2_8_32_58_inst0__clk = clk;

  assign ConfigRegister_2_8_32_58_inst0__config_addr[7:0] = config_config_addr[7:0];

  assign ConfigRegister_2_8_32_58_inst0__config_data[31:0] = config_config_data[31:0];

  assign ConfigRegister_2_8_32_58_inst0__config_en = config_write[0];

  assign ConfigRegister_2_8_32_58_inst0__reset = reset;

  assign MuxWrapper_4_1_inst15__S[1:0] = ConfigRegister_2_8_32_60_inst0__O[1:0];

  assign ZextWrapper_2_32_inst30__I[1:0] = ConfigRegister_2_8_32_60_inst0__O[1:0];

  assign ConfigRegister_2_8_32_60_inst0__clk = clk;

  assign ConfigRegister_2_8_32_60_inst0__config_addr[7:0] = config_config_addr[7:0];

  assign ConfigRegister_2_8_32_60_inst0__config_data[31:0] = config_config_data[31:0];

  assign ConfigRegister_2_8_32_60_inst0__config_en = config_write[0];

  assign ConfigRegister_2_8_32_60_inst0__reset = reset;

  assign MuxWrapper_4_1_inst16__S[1:0] = ConfigRegister_2_8_32_62_inst0__O[1:0];

  assign ZextWrapper_2_32_inst31__I[1:0] = ConfigRegister_2_8_32_62_inst0__O[1:0];

  assign ConfigRegister_2_8_32_62_inst0__clk = clk;

  assign ConfigRegister_2_8_32_62_inst0__config_addr[7:0] = config_config_addr[7:0];

  assign ConfigRegister_2_8_32_62_inst0__config_data[31:0] = config_config_data[31:0];

  assign ConfigRegister_2_8_32_62_inst0__config_en = config_write[0];

  assign ConfigRegister_2_8_32_62_inst0__reset = reset;

  assign MuxWrapper_4_1_inst17__S[1:0] = ConfigRegister_2_8_32_64_inst0__O[1:0];

  assign ZextWrapper_2_32_inst32__I[1:0] = ConfigRegister_2_8_32_64_inst0__O[1:0];

  assign ConfigRegister_2_8_32_64_inst0__clk = clk;

  assign ConfigRegister_2_8_32_64_inst0__config_addr[7:0] = config_config_addr[7:0];

  assign ConfigRegister_2_8_32_64_inst0__config_data[31:0] = config_config_data[31:0];

  assign ConfigRegister_2_8_32_64_inst0__config_en = config_write[0];

  assign ConfigRegister_2_8_32_64_inst0__reset = reset;

  assign MuxWrapper_4_1_inst18__S[1:0] = ConfigRegister_2_8_32_66_inst0__O[1:0];

  assign ZextWrapper_2_32_inst33__I[1:0] = ConfigRegister_2_8_32_66_inst0__O[1:0];

  assign ConfigRegister_2_8_32_66_inst0__clk = clk;

  assign ConfigRegister_2_8_32_66_inst0__config_addr[7:0] = config_config_addr[7:0];

  assign ConfigRegister_2_8_32_66_inst0__config_data[31:0] = config_config_data[31:0];

  assign ConfigRegister_2_8_32_66_inst0__config_en = config_write[0];

  assign ConfigRegister_2_8_32_66_inst0__reset = reset;

  assign MuxWrapper_4_1_inst19__S[1:0] = ConfigRegister_2_8_32_68_inst0__O[1:0];

  assign ZextWrapper_2_32_inst34__I[1:0] = ConfigRegister_2_8_32_68_inst0__O[1:0];

  assign ConfigRegister_2_8_32_68_inst0__clk = clk;

  assign ConfigRegister_2_8_32_68_inst0__config_addr[7:0] = config_config_addr[7:0];

  assign ConfigRegister_2_8_32_68_inst0__config_data[31:0] = config_config_data[31:0];

  assign ConfigRegister_2_8_32_68_inst0__config_en = config_write[0];

  assign ConfigRegister_2_8_32_68_inst0__reset = reset;

  assign MuxWrapper_4_1_inst3__S[1:0] = ConfigRegister_2_8_32_6_inst0__O[1:0];

  assign ZextWrapper_2_32_inst3__I[1:0] = ConfigRegister_2_8_32_6_inst0__O[1:0];

  assign ConfigRegister_2_8_32_6_inst0__clk = clk;

  assign ConfigRegister_2_8_32_6_inst0__config_addr[7:0] = config_config_addr[7:0];

  assign ConfigRegister_2_8_32_6_inst0__config_data[31:0] = config_config_data[31:0];

  assign ConfigRegister_2_8_32_6_inst0__config_en = config_write[0];

  assign ConfigRegister_2_8_32_6_inst0__reset = reset;

  assign MuxWrapper_4_16_inst15__S[1:0] = ConfigRegister_2_8_32_70_inst0__O[1:0];

  assign ZextWrapper_2_32_inst35__I[1:0] = ConfigRegister_2_8_32_70_inst0__O[1:0];

  assign ConfigRegister_2_8_32_70_inst0__clk = clk;

  assign ConfigRegister_2_8_32_70_inst0__config_addr[7:0] = config_config_addr[7:0];

  assign ConfigRegister_2_8_32_70_inst0__config_data[31:0] = config_config_data[31:0];

  assign ConfigRegister_2_8_32_70_inst0__config_en = config_write[0];

  assign ConfigRegister_2_8_32_70_inst0__reset = reset;

  assign MuxWrapper_4_16_inst16__S[1:0] = ConfigRegister_2_8_32_72_inst0__O[1:0];

  assign ZextWrapper_2_32_inst36__I[1:0] = ConfigRegister_2_8_32_72_inst0__O[1:0];

  assign ConfigRegister_2_8_32_72_inst0__clk = clk;

  assign ConfigRegister_2_8_32_72_inst0__config_addr[7:0] = config_config_addr[7:0];

  assign ConfigRegister_2_8_32_72_inst0__config_data[31:0] = config_config_data[31:0];

  assign ConfigRegister_2_8_32_72_inst0__config_en = config_write[0];

  assign ConfigRegister_2_8_32_72_inst0__reset = reset;

  assign MuxWrapper_4_16_inst17__S[1:0] = ConfigRegister_2_8_32_74_inst0__O[1:0];

  assign ZextWrapper_2_32_inst37__I[1:0] = ConfigRegister_2_8_32_74_inst0__O[1:0];

  assign ConfigRegister_2_8_32_74_inst0__clk = clk;

  assign ConfigRegister_2_8_32_74_inst0__config_addr[7:0] = config_config_addr[7:0];

  assign ConfigRegister_2_8_32_74_inst0__config_data[31:0] = config_config_data[31:0];

  assign ConfigRegister_2_8_32_74_inst0__config_en = config_write[0];

  assign ConfigRegister_2_8_32_74_inst0__reset = reset;

  assign MuxWrapper_4_16_inst18__S[1:0] = ConfigRegister_2_8_32_76_inst0__O[1:0];

  assign ZextWrapper_2_32_inst38__I[1:0] = ConfigRegister_2_8_32_76_inst0__O[1:0];

  assign ConfigRegister_2_8_32_76_inst0__clk = clk;

  assign ConfigRegister_2_8_32_76_inst0__config_addr[7:0] = config_config_addr[7:0];

  assign ConfigRegister_2_8_32_76_inst0__config_data[31:0] = config_config_data[31:0];

  assign ConfigRegister_2_8_32_76_inst0__config_en = config_write[0];

  assign ConfigRegister_2_8_32_76_inst0__reset = reset;

  assign MuxWrapper_4_16_inst19__S[1:0] = ConfigRegister_2_8_32_78_inst0__O[1:0];

  assign ZextWrapper_2_32_inst39__I[1:0] = ConfigRegister_2_8_32_78_inst0__O[1:0];

  assign ConfigRegister_2_8_32_78_inst0__clk = clk;

  assign ConfigRegister_2_8_32_78_inst0__config_addr[7:0] = config_config_addr[7:0];

  assign ConfigRegister_2_8_32_78_inst0__config_data[31:0] = config_config_data[31:0];

  assign ConfigRegister_2_8_32_78_inst0__config_en = config_write[0];

  assign ConfigRegister_2_8_32_78_inst0__reset = reset;

  assign MuxWrapper_4_1_inst4__S[1:0] = ConfigRegister_2_8_32_8_inst0__O[1:0];

  assign ZextWrapper_2_32_inst4__I[1:0] = ConfigRegister_2_8_32_8_inst0__O[1:0];

  assign ConfigRegister_2_8_32_8_inst0__clk = clk;

  assign ConfigRegister_2_8_32_8_inst0__config_addr[7:0] = config_config_addr[7:0];

  assign ConfigRegister_2_8_32_8_inst0__config_data[31:0] = config_config_data[31:0];

  assign ConfigRegister_2_8_32_8_inst0__config_en = config_write[0];

  assign ConfigRegister_2_8_32_8_inst0__reset = reset;

  assign MuxWrapper_2_16_inst0__I_0[15:0] = MuxWrapper_4_16_inst0__O[15:0];

  assign MuxWrapper_2_16_inst0__I_1[15:0] = reg_P_inst5__out[15:0];

  assign north_O_layer16_0[15:0] = MuxWrapper_2_16_inst0__O[15:0];

  assign MuxWrapper_2_16_inst1__I_0[15:0] = MuxWrapper_4_16_inst1__O[15:0];

  assign MuxWrapper_2_16_inst1__I_1[15:0] = reg_P_inst6__out[15:0];

  assign north_O_layer16_1[15:0] = MuxWrapper_2_16_inst1__O[15:0];

  assign MuxWrapper_2_16_inst10__I_0[15:0] = MuxWrapper_4_16_inst10__O[15:0];

  assign MuxWrapper_2_16_inst10__I_1[15:0] = reg_P_inst25__out[15:0];

  assign south_O_layer16_0[15:0] = MuxWrapper_2_16_inst10__O[15:0];

  assign MuxWrapper_2_16_inst11__I_0[15:0] = MuxWrapper_4_16_inst11__O[15:0];

  assign MuxWrapper_2_16_inst11__I_1[15:0] = reg_P_inst26__out[15:0];

  assign south_O_layer16_1[15:0] = MuxWrapper_2_16_inst11__O[15:0];

  assign MuxWrapper_2_16_inst12__I_0[15:0] = MuxWrapper_4_16_inst12__O[15:0];

  assign MuxWrapper_2_16_inst12__I_1[15:0] = reg_P_inst27__out[15:0];

  assign south_O_layer16_2[15:0] = MuxWrapper_2_16_inst12__O[15:0];

  assign MuxWrapper_2_16_inst13__I_0[15:0] = MuxWrapper_4_16_inst13__O[15:0];

  assign MuxWrapper_2_16_inst13__I_1[15:0] = reg_P_inst28__out[15:0];

  assign south_O_layer16_3[15:0] = MuxWrapper_2_16_inst13__O[15:0];

  assign MuxWrapper_2_16_inst14__I_0[15:0] = MuxWrapper_4_16_inst14__O[15:0];

  assign MuxWrapper_2_16_inst14__I_1[15:0] = reg_P_inst29__out[15:0];

  assign south_O_layer16_4[15:0] = MuxWrapper_2_16_inst14__O[15:0];

  assign MuxWrapper_2_16_inst15__I_0[15:0] = MuxWrapper_4_16_inst15__O[15:0];

  assign MuxWrapper_2_16_inst15__I_1[15:0] = reg_P_inst35__out[15:0];

  assign east_O_layer16_0[15:0] = MuxWrapper_2_16_inst15__O[15:0];

  assign MuxWrapper_2_16_inst16__I_0[15:0] = MuxWrapper_4_16_inst16__O[15:0];

  assign MuxWrapper_2_16_inst16__I_1[15:0] = reg_P_inst36__out[15:0];

  assign east_O_layer16_1[15:0] = MuxWrapper_2_16_inst16__O[15:0];

  assign MuxWrapper_2_16_inst17__I_0[15:0] = MuxWrapper_4_16_inst17__O[15:0];

  assign MuxWrapper_2_16_inst17__I_1[15:0] = reg_P_inst37__out[15:0];

  assign east_O_layer16_2[15:0] = MuxWrapper_2_16_inst17__O[15:0];

  assign MuxWrapper_2_16_inst18__I_0[15:0] = MuxWrapper_4_16_inst18__O[15:0];

  assign MuxWrapper_2_16_inst18__I_1[15:0] = reg_P_inst38__out[15:0];

  assign east_O_layer16_3[15:0] = MuxWrapper_2_16_inst18__O[15:0];

  assign MuxWrapper_2_16_inst19__I_0[15:0] = MuxWrapper_4_16_inst19__O[15:0];

  assign MuxWrapper_2_16_inst19__I_1[15:0] = reg_P_inst39__out[15:0];

  assign east_O_layer16_4[15:0] = MuxWrapper_2_16_inst19__O[15:0];

  assign MuxWrapper_2_16_inst2__I_0[15:0] = MuxWrapper_4_16_inst2__O[15:0];

  assign MuxWrapper_2_16_inst2__I_1[15:0] = reg_P_inst7__out[15:0];

  assign north_O_layer16_2[15:0] = MuxWrapper_2_16_inst2__O[15:0];

  assign MuxWrapper_2_16_inst3__I_0[15:0] = MuxWrapper_4_16_inst3__O[15:0];

  assign MuxWrapper_2_16_inst3__I_1[15:0] = reg_P_inst8__out[15:0];

  assign north_O_layer16_3[15:0] = MuxWrapper_2_16_inst3__O[15:0];

  assign MuxWrapper_2_16_inst4__I_0[15:0] = MuxWrapper_4_16_inst4__O[15:0];

  assign MuxWrapper_2_16_inst4__I_1[15:0] = reg_P_inst9__out[15:0];

  assign north_O_layer16_4[15:0] = MuxWrapper_2_16_inst4__O[15:0];

  assign MuxWrapper_2_16_inst5__I_0[15:0] = MuxWrapper_4_16_inst5__O[15:0];

  assign MuxWrapper_2_16_inst5__I_1[15:0] = reg_P_inst15__out[15:0];

  assign west_O_layer16_0[15:0] = MuxWrapper_2_16_inst5__O[15:0];

  assign MuxWrapper_2_16_inst6__I_0[15:0] = MuxWrapper_4_16_inst6__O[15:0];

  assign MuxWrapper_2_16_inst6__I_1[15:0] = reg_P_inst16__out[15:0];

  assign west_O_layer16_1[15:0] = MuxWrapper_2_16_inst6__O[15:0];

  assign MuxWrapper_2_16_inst7__I_0[15:0] = MuxWrapper_4_16_inst7__O[15:0];

  assign MuxWrapper_2_16_inst7__I_1[15:0] = reg_P_inst17__out[15:0];

  assign west_O_layer16_2[15:0] = MuxWrapper_2_16_inst7__O[15:0];

  assign MuxWrapper_2_16_inst8__I_0[15:0] = MuxWrapper_4_16_inst8__O[15:0];

  assign MuxWrapper_2_16_inst8__I_1[15:0] = reg_P_inst18__out[15:0];

  assign west_O_layer16_3[15:0] = MuxWrapper_2_16_inst8__O[15:0];

  assign MuxWrapper_2_16_inst9__I_0[15:0] = MuxWrapper_4_16_inst9__O[15:0];

  assign MuxWrapper_2_16_inst9__I_1[15:0] = reg_P_inst19__out[15:0];

  assign west_O_layer16_4[15:0] = MuxWrapper_2_16_inst9__O[15:0];

  assign MuxWrapper_2_1_inst0__I_0[0:0] = MuxWrapper_4_1_inst0__O[0:0];

  assign MuxWrapper_2_1_inst0__I_1[0:0] = reg_P_inst0__out[0:0];

  assign north_O_layer1_0[0:0] = MuxWrapper_2_1_inst0__O[0:0];

  assign MuxWrapper_2_1_inst1__I_0[0:0] = MuxWrapper_4_1_inst1__O[0:0];

  assign MuxWrapper_2_1_inst1__I_1[0:0] = reg_P_inst1__out[0:0];

  assign north_O_layer1_1[0:0] = MuxWrapper_2_1_inst1__O[0:0];

  assign MuxWrapper_2_1_inst10__I_0[0:0] = MuxWrapper_4_1_inst10__O[0:0];

  assign MuxWrapper_2_1_inst10__I_1[0:0] = reg_P_inst20__out[0:0];

  assign south_O_layer1_0[0:0] = MuxWrapper_2_1_inst10__O[0:0];

  assign MuxWrapper_2_1_inst11__I_0[0:0] = MuxWrapper_4_1_inst11__O[0:0];

  assign MuxWrapper_2_1_inst11__I_1[0:0] = reg_P_inst21__out[0:0];

  assign south_O_layer1_1[0:0] = MuxWrapper_2_1_inst11__O[0:0];

  assign MuxWrapper_2_1_inst12__I_0[0:0] = MuxWrapper_4_1_inst12__O[0:0];

  assign MuxWrapper_2_1_inst12__I_1[0:0] = reg_P_inst22__out[0:0];

  assign south_O_layer1_2[0:0] = MuxWrapper_2_1_inst12__O[0:0];

  assign MuxWrapper_2_1_inst13__I_0[0:0] = MuxWrapper_4_1_inst13__O[0:0];

  assign MuxWrapper_2_1_inst13__I_1[0:0] = reg_P_inst23__out[0:0];

  assign south_O_layer1_3[0:0] = MuxWrapper_2_1_inst13__O[0:0];

  assign MuxWrapper_2_1_inst14__I_0[0:0] = MuxWrapper_4_1_inst14__O[0:0];

  assign MuxWrapper_2_1_inst14__I_1[0:0] = reg_P_inst24__out[0:0];

  assign south_O_layer1_4[0:0] = MuxWrapper_2_1_inst14__O[0:0];

  assign MuxWrapper_2_1_inst15__I_0[0:0] = MuxWrapper_4_1_inst15__O[0:0];

  assign MuxWrapper_2_1_inst15__I_1[0:0] = reg_P_inst30__out[0:0];

  assign east_O_layer1_0[0:0] = MuxWrapper_2_1_inst15__O[0:0];

  assign MuxWrapper_2_1_inst16__I_0[0:0] = MuxWrapper_4_1_inst16__O[0:0];

  assign MuxWrapper_2_1_inst16__I_1[0:0] = reg_P_inst31__out[0:0];

  assign east_O_layer1_1[0:0] = MuxWrapper_2_1_inst16__O[0:0];

  assign MuxWrapper_2_1_inst17__I_0[0:0] = MuxWrapper_4_1_inst17__O[0:0];

  assign MuxWrapper_2_1_inst17__I_1[0:0] = reg_P_inst32__out[0:0];

  assign east_O_layer1_2[0:0] = MuxWrapper_2_1_inst17__O[0:0];

  assign MuxWrapper_2_1_inst18__I_0[0:0] = MuxWrapper_4_1_inst18__O[0:0];

  assign MuxWrapper_2_1_inst18__I_1[0:0] = reg_P_inst33__out[0:0];

  assign east_O_layer1_3[0:0] = MuxWrapper_2_1_inst18__O[0:0];

  assign MuxWrapper_2_1_inst19__I_0[0:0] = MuxWrapper_4_1_inst19__O[0:0];

  assign MuxWrapper_2_1_inst19__I_1[0:0] = reg_P_inst34__out[0:0];

  assign east_O_layer1_4[0:0] = MuxWrapper_2_1_inst19__O[0:0];

  assign MuxWrapper_2_1_inst2__I_0[0:0] = MuxWrapper_4_1_inst2__O[0:0];

  assign MuxWrapper_2_1_inst2__I_1[0:0] = reg_P_inst2__out[0:0];

  assign north_O_layer1_2[0:0] = MuxWrapper_2_1_inst2__O[0:0];

  assign MuxWrapper_2_1_inst3__I_0[0:0] = MuxWrapper_4_1_inst3__O[0:0];

  assign MuxWrapper_2_1_inst3__I_1[0:0] = reg_P_inst3__out[0:0];

  assign north_O_layer1_3[0:0] = MuxWrapper_2_1_inst3__O[0:0];

  assign MuxWrapper_2_1_inst4__I_0[0:0] = MuxWrapper_4_1_inst4__O[0:0];

  assign MuxWrapper_2_1_inst4__I_1[0:0] = reg_P_inst4__out[0:0];

  assign north_O_layer1_4[0:0] = MuxWrapper_2_1_inst4__O[0:0];

  assign MuxWrapper_2_1_inst5__I_0[0:0] = MuxWrapper_4_1_inst5__O[0:0];

  assign MuxWrapper_2_1_inst5__I_1[0:0] = reg_P_inst10__out[0:0];

  assign west_O_layer1_0[0:0] = MuxWrapper_2_1_inst5__O[0:0];

  assign MuxWrapper_2_1_inst6__I_0[0:0] = MuxWrapper_4_1_inst6__O[0:0];

  assign MuxWrapper_2_1_inst6__I_1[0:0] = reg_P_inst11__out[0:0];

  assign west_O_layer1_1[0:0] = MuxWrapper_2_1_inst6__O[0:0];

  assign MuxWrapper_2_1_inst7__I_0[0:0] = MuxWrapper_4_1_inst7__O[0:0];

  assign MuxWrapper_2_1_inst7__I_1[0:0] = reg_P_inst12__out[0:0];

  assign west_O_layer1_2[0:0] = MuxWrapper_2_1_inst7__O[0:0];

  assign MuxWrapper_2_1_inst8__I_0[0:0] = MuxWrapper_4_1_inst8__O[0:0];

  assign MuxWrapper_2_1_inst8__I_1[0:0] = reg_P_inst13__out[0:0];

  assign west_O_layer1_3[0:0] = MuxWrapper_2_1_inst8__O[0:0];

  assign MuxWrapper_2_1_inst9__I_0[0:0] = MuxWrapper_4_1_inst9__O[0:0];

  assign MuxWrapper_2_1_inst9__I_1[0:0] = reg_P_inst14__out[0:0];

  assign west_O_layer1_4[0:0] = MuxWrapper_2_1_inst9__O[0:0];

  assign MuxWrapper_4_16_inst0__I_0[15:0] = west_I_layer16_0[15:0];

  assign MuxWrapper_4_16_inst0__I_1[15:0] = south_I_layer16_0[15:0];

  assign MuxWrapper_4_16_inst0__I_2[15:0] = east_I_layer16_0[15:0];

  assign MuxWrapper_4_16_inst0__I_3[15:0] = res[15:0];

  assign reg_P_inst5__in[15:0] = MuxWrapper_4_16_inst0__O[15:0];

  assign MuxWrapper_4_16_inst1__I_0[15:0] = west_I_layer16_1[15:0];

  assign MuxWrapper_4_16_inst1__I_1[15:0] = south_I_layer16_1[15:0];

  assign MuxWrapper_4_16_inst1__I_2[15:0] = east_I_layer16_1[15:0];

  assign MuxWrapper_4_16_inst1__I_3[15:0] = res[15:0];

  assign reg_P_inst6__in[15:0] = MuxWrapper_4_16_inst1__O[15:0];

  assign MuxWrapper_4_16_inst10__I_0[15:0] = north_I_layer16_0[15:0];

  assign MuxWrapper_4_16_inst10__I_1[15:0] = west_I_layer16_0[15:0];

  assign MuxWrapper_4_16_inst10__I_2[15:0] = east_I_layer16_0[15:0];

  assign MuxWrapper_4_16_inst10__I_3[15:0] = res[15:0];

  assign reg_P_inst25__in[15:0] = MuxWrapper_4_16_inst10__O[15:0];

  assign MuxWrapper_4_16_inst11__I_0[15:0] = north_I_layer16_1[15:0];

  assign MuxWrapper_4_16_inst11__I_1[15:0] = west_I_layer16_1[15:0];

  assign MuxWrapper_4_16_inst11__I_2[15:0] = east_I_layer16_1[15:0];

  assign MuxWrapper_4_16_inst11__I_3[15:0] = res[15:0];

  assign reg_P_inst26__in[15:0] = MuxWrapper_4_16_inst11__O[15:0];

  assign MuxWrapper_4_16_inst12__I_0[15:0] = north_I_layer16_2[15:0];

  assign MuxWrapper_4_16_inst12__I_1[15:0] = west_I_layer16_2[15:0];

  assign MuxWrapper_4_16_inst12__I_2[15:0] = east_I_layer16_2[15:0];

  assign MuxWrapper_4_16_inst12__I_3[15:0] = res[15:0];

  assign reg_P_inst27__in[15:0] = MuxWrapper_4_16_inst12__O[15:0];

  assign MuxWrapper_4_16_inst13__I_0[15:0] = north_I_layer16_3[15:0];

  assign MuxWrapper_4_16_inst13__I_1[15:0] = west_I_layer16_3[15:0];

  assign MuxWrapper_4_16_inst13__I_2[15:0] = east_I_layer16_3[15:0];

  assign MuxWrapper_4_16_inst13__I_3[15:0] = res[15:0];

  assign reg_P_inst28__in[15:0] = MuxWrapper_4_16_inst13__O[15:0];

  assign MuxWrapper_4_16_inst14__I_0[15:0] = north_I_layer16_4[15:0];

  assign MuxWrapper_4_16_inst14__I_1[15:0] = west_I_layer16_4[15:0];

  assign MuxWrapper_4_16_inst14__I_2[15:0] = east_I_layer16_4[15:0];

  assign MuxWrapper_4_16_inst14__I_3[15:0] = res[15:0];

  assign reg_P_inst29__in[15:0] = MuxWrapper_4_16_inst14__O[15:0];

  assign MuxWrapper_4_16_inst15__I_0[15:0] = north_I_layer16_0[15:0];

  assign MuxWrapper_4_16_inst15__I_1[15:0] = west_I_layer16_0[15:0];

  assign MuxWrapper_4_16_inst15__I_2[15:0] = south_I_layer16_0[15:0];

  assign MuxWrapper_4_16_inst15__I_3[15:0] = res[15:0];

  assign reg_P_inst35__in[15:0] = MuxWrapper_4_16_inst15__O[15:0];

  assign MuxWrapper_4_16_inst16__I_0[15:0] = north_I_layer16_1[15:0];

  assign MuxWrapper_4_16_inst16__I_1[15:0] = west_I_layer16_1[15:0];

  assign MuxWrapper_4_16_inst16__I_2[15:0] = south_I_layer16_1[15:0];

  assign MuxWrapper_4_16_inst16__I_3[15:0] = res[15:0];

  assign reg_P_inst36__in[15:0] = MuxWrapper_4_16_inst16__O[15:0];

  assign MuxWrapper_4_16_inst17__I_0[15:0] = north_I_layer16_2[15:0];

  assign MuxWrapper_4_16_inst17__I_1[15:0] = west_I_layer16_2[15:0];

  assign MuxWrapper_4_16_inst17__I_2[15:0] = south_I_layer16_2[15:0];

  assign MuxWrapper_4_16_inst17__I_3[15:0] = res[15:0];

  assign reg_P_inst37__in[15:0] = MuxWrapper_4_16_inst17__O[15:0];

  assign MuxWrapper_4_16_inst18__I_0[15:0] = north_I_layer16_3[15:0];

  assign MuxWrapper_4_16_inst18__I_1[15:0] = west_I_layer16_3[15:0];

  assign MuxWrapper_4_16_inst18__I_2[15:0] = south_I_layer16_3[15:0];

  assign MuxWrapper_4_16_inst18__I_3[15:0] = res[15:0];

  assign reg_P_inst38__in[15:0] = MuxWrapper_4_16_inst18__O[15:0];

  assign MuxWrapper_4_16_inst19__I_0[15:0] = north_I_layer16_4[15:0];

  assign MuxWrapper_4_16_inst19__I_1[15:0] = west_I_layer16_4[15:0];

  assign MuxWrapper_4_16_inst19__I_2[15:0] = south_I_layer16_4[15:0];

  assign MuxWrapper_4_16_inst19__I_3[15:0] = res[15:0];

  assign reg_P_inst39__in[15:0] = MuxWrapper_4_16_inst19__O[15:0];

  assign MuxWrapper_4_16_inst2__I_0[15:0] = west_I_layer16_2[15:0];

  assign MuxWrapper_4_16_inst2__I_1[15:0] = south_I_layer16_2[15:0];

  assign MuxWrapper_4_16_inst2__I_2[15:0] = east_I_layer16_2[15:0];

  assign MuxWrapper_4_16_inst2__I_3[15:0] = res[15:0];

  assign reg_P_inst7__in[15:0] = MuxWrapper_4_16_inst2__O[15:0];

  assign MuxWrapper_4_16_inst3__I_0[15:0] = west_I_layer16_3[15:0];

  assign MuxWrapper_4_16_inst3__I_1[15:0] = south_I_layer16_3[15:0];

  assign MuxWrapper_4_16_inst3__I_2[15:0] = east_I_layer16_3[15:0];

  assign MuxWrapper_4_16_inst3__I_3[15:0] = res[15:0];

  assign reg_P_inst8__in[15:0] = MuxWrapper_4_16_inst3__O[15:0];

  assign MuxWrapper_4_16_inst4__I_0[15:0] = west_I_layer16_4[15:0];

  assign MuxWrapper_4_16_inst4__I_1[15:0] = south_I_layer16_4[15:0];

  assign MuxWrapper_4_16_inst4__I_2[15:0] = east_I_layer16_4[15:0];

  assign MuxWrapper_4_16_inst4__I_3[15:0] = res[15:0];

  assign reg_P_inst9__in[15:0] = MuxWrapper_4_16_inst4__O[15:0];

  assign MuxWrapper_4_16_inst5__I_0[15:0] = north_I_layer16_0[15:0];

  assign MuxWrapper_4_16_inst5__I_1[15:0] = south_I_layer16_0[15:0];

  assign MuxWrapper_4_16_inst5__I_2[15:0] = east_I_layer16_0[15:0];

  assign MuxWrapper_4_16_inst5__I_3[15:0] = res[15:0];

  assign reg_P_inst15__in[15:0] = MuxWrapper_4_16_inst5__O[15:0];

  assign MuxWrapper_4_16_inst6__I_0[15:0] = north_I_layer16_1[15:0];

  assign MuxWrapper_4_16_inst6__I_1[15:0] = south_I_layer16_1[15:0];

  assign MuxWrapper_4_16_inst6__I_2[15:0] = east_I_layer16_1[15:0];

  assign MuxWrapper_4_16_inst6__I_3[15:0] = res[15:0];

  assign reg_P_inst16__in[15:0] = MuxWrapper_4_16_inst6__O[15:0];

  assign MuxWrapper_4_16_inst7__I_0[15:0] = north_I_layer16_2[15:0];

  assign MuxWrapper_4_16_inst7__I_1[15:0] = south_I_layer16_2[15:0];

  assign MuxWrapper_4_16_inst7__I_2[15:0] = east_I_layer16_2[15:0];

  assign MuxWrapper_4_16_inst7__I_3[15:0] = res[15:0];

  assign reg_P_inst17__in[15:0] = MuxWrapper_4_16_inst7__O[15:0];

  assign MuxWrapper_4_16_inst8__I_0[15:0] = north_I_layer16_3[15:0];

  assign MuxWrapper_4_16_inst8__I_1[15:0] = south_I_layer16_3[15:0];

  assign MuxWrapper_4_16_inst8__I_2[15:0] = east_I_layer16_3[15:0];

  assign MuxWrapper_4_16_inst8__I_3[15:0] = res[15:0];

  assign reg_P_inst18__in[15:0] = MuxWrapper_4_16_inst8__O[15:0];

  assign MuxWrapper_4_16_inst9__I_0[15:0] = north_I_layer16_4[15:0];

  assign MuxWrapper_4_16_inst9__I_1[15:0] = south_I_layer16_4[15:0];

  assign MuxWrapper_4_16_inst9__I_2[15:0] = east_I_layer16_4[15:0];

  assign MuxWrapper_4_16_inst9__I_3[15:0] = res[15:0];

  assign reg_P_inst19__in[15:0] = MuxWrapper_4_16_inst9__O[15:0];

  assign MuxWrapper_4_1_inst0__I_0[0:0] = west_I_layer1_0[0:0];

  assign MuxWrapper_4_1_inst0__I_1[0:0] = south_I_layer1_0[0:0];

  assign MuxWrapper_4_1_inst0__I_2[0:0] = east_I_layer1_0[0:0];

  assign MuxWrapper_4_1_inst0__I_3[0:0] = res_p[0:0];

  assign reg_P_inst0__in[0:0] = MuxWrapper_4_1_inst0__O[0:0];

  assign MuxWrapper_4_1_inst1__I_0[0:0] = west_I_layer1_1[0:0];

  assign MuxWrapper_4_1_inst1__I_1[0:0] = south_I_layer1_1[0:0];

  assign MuxWrapper_4_1_inst1__I_2[0:0] = east_I_layer1_1[0:0];

  assign MuxWrapper_4_1_inst1__I_3[0:0] = res_p[0:0];

  assign reg_P_inst1__in[0:0] = MuxWrapper_4_1_inst1__O[0:0];

  assign MuxWrapper_4_1_inst10__I_0[0:0] = north_I_layer1_0[0:0];

  assign MuxWrapper_4_1_inst10__I_1[0:0] = west_I_layer1_0[0:0];

  assign MuxWrapper_4_1_inst10__I_2[0:0] = east_I_layer1_0[0:0];

  assign MuxWrapper_4_1_inst10__I_3[0:0] = res_p[0:0];

  assign reg_P_inst20__in[0:0] = MuxWrapper_4_1_inst10__O[0:0];

  assign MuxWrapper_4_1_inst11__I_0[0:0] = north_I_layer1_1[0:0];

  assign MuxWrapper_4_1_inst11__I_1[0:0] = west_I_layer1_1[0:0];

  assign MuxWrapper_4_1_inst11__I_2[0:0] = east_I_layer1_1[0:0];

  assign MuxWrapper_4_1_inst11__I_3[0:0] = res_p[0:0];

  assign reg_P_inst21__in[0:0] = MuxWrapper_4_1_inst11__O[0:0];

  assign MuxWrapper_4_1_inst12__I_0[0:0] = north_I_layer1_2[0:0];

  assign MuxWrapper_4_1_inst12__I_1[0:0] = west_I_layer1_2[0:0];

  assign MuxWrapper_4_1_inst12__I_2[0:0] = east_I_layer1_2[0:0];

  assign MuxWrapper_4_1_inst12__I_3[0:0] = res_p[0:0];

  assign reg_P_inst22__in[0:0] = MuxWrapper_4_1_inst12__O[0:0];

  assign MuxWrapper_4_1_inst13__I_0[0:0] = north_I_layer1_3[0:0];

  assign MuxWrapper_4_1_inst13__I_1[0:0] = west_I_layer1_3[0:0];

  assign MuxWrapper_4_1_inst13__I_2[0:0] = east_I_layer1_3[0:0];

  assign MuxWrapper_4_1_inst13__I_3[0:0] = res_p[0:0];

  assign reg_P_inst23__in[0:0] = MuxWrapper_4_1_inst13__O[0:0];

  assign MuxWrapper_4_1_inst14__I_0[0:0] = north_I_layer1_4[0:0];

  assign MuxWrapper_4_1_inst14__I_1[0:0] = west_I_layer1_4[0:0];

  assign MuxWrapper_4_1_inst14__I_2[0:0] = east_I_layer1_4[0:0];

  assign MuxWrapper_4_1_inst14__I_3[0:0] = res_p[0:0];

  assign reg_P_inst24__in[0:0] = MuxWrapper_4_1_inst14__O[0:0];

  assign MuxWrapper_4_1_inst15__I_0[0:0] = north_I_layer1_0[0:0];

  assign MuxWrapper_4_1_inst15__I_1[0:0] = west_I_layer1_0[0:0];

  assign MuxWrapper_4_1_inst15__I_2[0:0] = south_I_layer1_0[0:0];

  assign MuxWrapper_4_1_inst15__I_3[0:0] = res_p[0:0];

  assign reg_P_inst30__in[0:0] = MuxWrapper_4_1_inst15__O[0:0];

  assign MuxWrapper_4_1_inst16__I_0[0:0] = north_I_layer1_1[0:0];

  assign MuxWrapper_4_1_inst16__I_1[0:0] = west_I_layer1_1[0:0];

  assign MuxWrapper_4_1_inst16__I_2[0:0] = south_I_layer1_1[0:0];

  assign MuxWrapper_4_1_inst16__I_3[0:0] = res_p[0:0];

  assign reg_P_inst31__in[0:0] = MuxWrapper_4_1_inst16__O[0:0];

  assign MuxWrapper_4_1_inst17__I_0[0:0] = north_I_layer1_2[0:0];

  assign MuxWrapper_4_1_inst17__I_1[0:0] = west_I_layer1_2[0:0];

  assign MuxWrapper_4_1_inst17__I_2[0:0] = south_I_layer1_2[0:0];

  assign MuxWrapper_4_1_inst17__I_3[0:0] = res_p[0:0];

  assign reg_P_inst32__in[0:0] = MuxWrapper_4_1_inst17__O[0:0];

  assign MuxWrapper_4_1_inst18__I_0[0:0] = north_I_layer1_3[0:0];

  assign MuxWrapper_4_1_inst18__I_1[0:0] = west_I_layer1_3[0:0];

  assign MuxWrapper_4_1_inst18__I_2[0:0] = south_I_layer1_3[0:0];

  assign MuxWrapper_4_1_inst18__I_3[0:0] = res_p[0:0];

  assign reg_P_inst33__in[0:0] = MuxWrapper_4_1_inst18__O[0:0];

  assign MuxWrapper_4_1_inst19__I_0[0:0] = north_I_layer1_4[0:0];

  assign MuxWrapper_4_1_inst19__I_1[0:0] = west_I_layer1_4[0:0];

  assign MuxWrapper_4_1_inst19__I_2[0:0] = south_I_layer1_4[0:0];

  assign MuxWrapper_4_1_inst19__I_3[0:0] = res_p[0:0];

  assign reg_P_inst34__in[0:0] = MuxWrapper_4_1_inst19__O[0:0];

  assign MuxWrapper_4_1_inst2__I_0[0:0] = west_I_layer1_2[0:0];

  assign MuxWrapper_4_1_inst2__I_1[0:0] = south_I_layer1_2[0:0];

  assign MuxWrapper_4_1_inst2__I_2[0:0] = east_I_layer1_2[0:0];

  assign MuxWrapper_4_1_inst2__I_3[0:0] = res_p[0:0];

  assign reg_P_inst2__in[0:0] = MuxWrapper_4_1_inst2__O[0:0];

  assign MuxWrapper_4_1_inst3__I_0[0:0] = west_I_layer1_3[0:0];

  assign MuxWrapper_4_1_inst3__I_1[0:0] = south_I_layer1_3[0:0];

  assign MuxWrapper_4_1_inst3__I_2[0:0] = east_I_layer1_3[0:0];

  assign MuxWrapper_4_1_inst3__I_3[0:0] = res_p[0:0];

  assign reg_P_inst3__in[0:0] = MuxWrapper_4_1_inst3__O[0:0];

  assign MuxWrapper_4_1_inst4__I_0[0:0] = west_I_layer1_4[0:0];

  assign MuxWrapper_4_1_inst4__I_1[0:0] = south_I_layer1_4[0:0];

  assign MuxWrapper_4_1_inst4__I_2[0:0] = east_I_layer1_4[0:0];

  assign MuxWrapper_4_1_inst4__I_3[0:0] = res_p[0:0];

  assign reg_P_inst4__in[0:0] = MuxWrapper_4_1_inst4__O[0:0];

  assign MuxWrapper_4_1_inst5__I_0[0:0] = north_I_layer1_0[0:0];

  assign MuxWrapper_4_1_inst5__I_1[0:0] = south_I_layer1_0[0:0];

  assign MuxWrapper_4_1_inst5__I_2[0:0] = east_I_layer1_0[0:0];

  assign MuxWrapper_4_1_inst5__I_3[0:0] = res_p[0:0];

  assign reg_P_inst10__in[0:0] = MuxWrapper_4_1_inst5__O[0:0];

  assign MuxWrapper_4_1_inst6__I_0[0:0] = north_I_layer1_1[0:0];

  assign MuxWrapper_4_1_inst6__I_1[0:0] = south_I_layer1_1[0:0];

  assign MuxWrapper_4_1_inst6__I_2[0:0] = east_I_layer1_1[0:0];

  assign MuxWrapper_4_1_inst6__I_3[0:0] = res_p[0:0];

  assign reg_P_inst11__in[0:0] = MuxWrapper_4_1_inst6__O[0:0];

  assign MuxWrapper_4_1_inst7__I_0[0:0] = north_I_layer1_2[0:0];

  assign MuxWrapper_4_1_inst7__I_1[0:0] = south_I_layer1_2[0:0];

  assign MuxWrapper_4_1_inst7__I_2[0:0] = east_I_layer1_2[0:0];

  assign MuxWrapper_4_1_inst7__I_3[0:0] = res_p[0:0];

  assign reg_P_inst12__in[0:0] = MuxWrapper_4_1_inst7__O[0:0];

  assign MuxWrapper_4_1_inst8__I_0[0:0] = north_I_layer1_3[0:0];

  assign MuxWrapper_4_1_inst8__I_1[0:0] = south_I_layer1_3[0:0];

  assign MuxWrapper_4_1_inst8__I_2[0:0] = east_I_layer1_3[0:0];

  assign MuxWrapper_4_1_inst8__I_3[0:0] = res_p[0:0];

  assign reg_P_inst13__in[0:0] = MuxWrapper_4_1_inst8__O[0:0];

  assign MuxWrapper_4_1_inst9__I_0[0:0] = north_I_layer1_4[0:0];

  assign MuxWrapper_4_1_inst9__I_1[0:0] = south_I_layer1_4[0:0];

  assign MuxWrapper_4_1_inst9__I_2[0:0] = east_I_layer1_4[0:0];

  assign MuxWrapper_4_1_inst9__I_3[0:0] = res_p[0:0];

  assign reg_P_inst14__in[0:0] = MuxWrapper_4_1_inst9__O[0:0];

  assign MuxWrapper_80_32_inst0__I_0[31:0] = ZextWrapper_2_32_inst0__O[31:0];

  assign MuxWrapper_80_32_inst0__I_1[31:0] = ZextWrapper_1_32_inst0__O[31:0];

  assign MuxWrapper_80_32_inst0__I_10[31:0] = ZextWrapper_2_32_inst5__O[31:0];

  assign MuxWrapper_80_32_inst0__I_11[31:0] = ZextWrapper_1_32_inst5__O[31:0];

  assign MuxWrapper_80_32_inst0__I_12[31:0] = ZextWrapper_2_32_inst6__O[31:0];

  assign MuxWrapper_80_32_inst0__I_13[31:0] = ZextWrapper_1_32_inst6__O[31:0];

  assign MuxWrapper_80_32_inst0__I_14[31:0] = ZextWrapper_2_32_inst7__O[31:0];

  assign MuxWrapper_80_32_inst0__I_15[31:0] = ZextWrapper_1_32_inst7__O[31:0];

  assign MuxWrapper_80_32_inst0__I_16[31:0] = ZextWrapper_2_32_inst8__O[31:0];

  assign MuxWrapper_80_32_inst0__I_17[31:0] = ZextWrapper_1_32_inst8__O[31:0];

  assign MuxWrapper_80_32_inst0__I_18[31:0] = ZextWrapper_2_32_inst9__O[31:0];

  assign MuxWrapper_80_32_inst0__I_19[31:0] = ZextWrapper_1_32_inst9__O[31:0];

  assign MuxWrapper_80_32_inst0__I_2[31:0] = ZextWrapper_2_32_inst1__O[31:0];

  assign MuxWrapper_80_32_inst0__I_20[31:0] = ZextWrapper_2_32_inst10__O[31:0];

  assign MuxWrapper_80_32_inst0__I_21[31:0] = ZextWrapper_1_32_inst10__O[31:0];

  assign MuxWrapper_80_32_inst0__I_22[31:0] = ZextWrapper_2_32_inst11__O[31:0];

  assign MuxWrapper_80_32_inst0__I_23[31:0] = ZextWrapper_1_32_inst11__O[31:0];

  assign MuxWrapper_80_32_inst0__I_24[31:0] = ZextWrapper_2_32_inst12__O[31:0];

  assign MuxWrapper_80_32_inst0__I_25[31:0] = ZextWrapper_1_32_inst12__O[31:0];

  assign MuxWrapper_80_32_inst0__I_26[31:0] = ZextWrapper_2_32_inst13__O[31:0];

  assign MuxWrapper_80_32_inst0__I_27[31:0] = ZextWrapper_1_32_inst13__O[31:0];

  assign MuxWrapper_80_32_inst0__I_28[31:0] = ZextWrapper_2_32_inst14__O[31:0];

  assign MuxWrapper_80_32_inst0__I_29[31:0] = ZextWrapper_1_32_inst14__O[31:0];

  assign MuxWrapper_80_32_inst0__I_3[31:0] = ZextWrapper_1_32_inst1__O[31:0];

  assign MuxWrapper_80_32_inst0__I_30[31:0] = ZextWrapper_2_32_inst15__O[31:0];

  assign MuxWrapper_80_32_inst0__I_31[31:0] = ZextWrapper_1_32_inst15__O[31:0];

  assign MuxWrapper_80_32_inst0__I_32[31:0] = ZextWrapper_2_32_inst16__O[31:0];

  assign MuxWrapper_80_32_inst0__I_33[31:0] = ZextWrapper_1_32_inst16__O[31:0];

  assign MuxWrapper_80_32_inst0__I_34[31:0] = ZextWrapper_2_32_inst17__O[31:0];

  assign MuxWrapper_80_32_inst0__I_35[31:0] = ZextWrapper_1_32_inst17__O[31:0];

  assign MuxWrapper_80_32_inst0__I_36[31:0] = ZextWrapper_2_32_inst18__O[31:0];

  assign MuxWrapper_80_32_inst0__I_37[31:0] = ZextWrapper_1_32_inst18__O[31:0];

  assign MuxWrapper_80_32_inst0__I_38[31:0] = ZextWrapper_2_32_inst19__O[31:0];

  assign MuxWrapper_80_32_inst0__I_39[31:0] = ZextWrapper_1_32_inst19__O[31:0];

  assign MuxWrapper_80_32_inst0__I_4[31:0] = ZextWrapper_2_32_inst2__O[31:0];

  assign MuxWrapper_80_32_inst0__I_40[31:0] = ZextWrapper_2_32_inst20__O[31:0];

  assign MuxWrapper_80_32_inst0__I_41[31:0] = ZextWrapper_1_32_inst20__O[31:0];

  assign MuxWrapper_80_32_inst0__I_42[31:0] = ZextWrapper_2_32_inst21__O[31:0];

  assign MuxWrapper_80_32_inst0__I_43[31:0] = ZextWrapper_1_32_inst21__O[31:0];

  assign MuxWrapper_80_32_inst0__I_44[31:0] = ZextWrapper_2_32_inst22__O[31:0];

  assign MuxWrapper_80_32_inst0__I_45[31:0] = ZextWrapper_1_32_inst22__O[31:0];

  assign MuxWrapper_80_32_inst0__I_46[31:0] = ZextWrapper_2_32_inst23__O[31:0];

  assign MuxWrapper_80_32_inst0__I_47[31:0] = ZextWrapper_1_32_inst23__O[31:0];

  assign MuxWrapper_80_32_inst0__I_48[31:0] = ZextWrapper_2_32_inst24__O[31:0];

  assign MuxWrapper_80_32_inst0__I_49[31:0] = ZextWrapper_1_32_inst24__O[31:0];

  assign MuxWrapper_80_32_inst0__I_5[31:0] = ZextWrapper_1_32_inst2__O[31:0];

  assign MuxWrapper_80_32_inst0__I_50[31:0] = ZextWrapper_2_32_inst25__O[31:0];

  assign MuxWrapper_80_32_inst0__I_51[31:0] = ZextWrapper_1_32_inst25__O[31:0];

  assign MuxWrapper_80_32_inst0__I_52[31:0] = ZextWrapper_2_32_inst26__O[31:0];

  assign MuxWrapper_80_32_inst0__I_53[31:0] = ZextWrapper_1_32_inst26__O[31:0];

  assign MuxWrapper_80_32_inst0__I_54[31:0] = ZextWrapper_2_32_inst27__O[31:0];

  assign MuxWrapper_80_32_inst0__I_55[31:0] = ZextWrapper_1_32_inst27__O[31:0];

  assign MuxWrapper_80_32_inst0__I_56[31:0] = ZextWrapper_2_32_inst28__O[31:0];

  assign MuxWrapper_80_32_inst0__I_57[31:0] = ZextWrapper_1_32_inst28__O[31:0];

  assign MuxWrapper_80_32_inst0__I_58[31:0] = ZextWrapper_2_32_inst29__O[31:0];

  assign MuxWrapper_80_32_inst0__I_59[31:0] = ZextWrapper_1_32_inst29__O[31:0];

  assign MuxWrapper_80_32_inst0__I_6[31:0] = ZextWrapper_2_32_inst3__O[31:0];

  assign MuxWrapper_80_32_inst0__I_60[31:0] = ZextWrapper_2_32_inst30__O[31:0];

  assign MuxWrapper_80_32_inst0__I_61[31:0] = ZextWrapper_1_32_inst30__O[31:0];

  assign MuxWrapper_80_32_inst0__I_62[31:0] = ZextWrapper_2_32_inst31__O[31:0];

  assign MuxWrapper_80_32_inst0__I_63[31:0] = ZextWrapper_1_32_inst31__O[31:0];

  assign MuxWrapper_80_32_inst0__I_64[31:0] = ZextWrapper_2_32_inst32__O[31:0];

  assign MuxWrapper_80_32_inst0__I_65[31:0] = ZextWrapper_1_32_inst32__O[31:0];

  assign MuxWrapper_80_32_inst0__I_66[31:0] = ZextWrapper_2_32_inst33__O[31:0];

  assign MuxWrapper_80_32_inst0__I_67[31:0] = ZextWrapper_1_32_inst33__O[31:0];

  assign MuxWrapper_80_32_inst0__I_68[31:0] = ZextWrapper_2_32_inst34__O[31:0];

  assign MuxWrapper_80_32_inst0__I_69[31:0] = ZextWrapper_1_32_inst34__O[31:0];

  assign MuxWrapper_80_32_inst0__I_7[31:0] = ZextWrapper_1_32_inst3__O[31:0];

  assign MuxWrapper_80_32_inst0__I_70[31:0] = ZextWrapper_2_32_inst35__O[31:0];

  assign MuxWrapper_80_32_inst0__I_71[31:0] = ZextWrapper_1_32_inst35__O[31:0];

  assign MuxWrapper_80_32_inst0__I_72[31:0] = ZextWrapper_2_32_inst36__O[31:0];

  assign MuxWrapper_80_32_inst0__I_73[31:0] = ZextWrapper_1_32_inst36__O[31:0];

  assign MuxWrapper_80_32_inst0__I_74[31:0] = ZextWrapper_2_32_inst37__O[31:0];

  assign MuxWrapper_80_32_inst0__I_75[31:0] = ZextWrapper_1_32_inst37__O[31:0];

  assign MuxWrapper_80_32_inst0__I_76[31:0] = ZextWrapper_2_32_inst38__O[31:0];

  assign MuxWrapper_80_32_inst0__I_77[31:0] = ZextWrapper_1_32_inst38__O[31:0];

  assign MuxWrapper_80_32_inst0__I_78[31:0] = ZextWrapper_2_32_inst39__O[31:0];

  assign MuxWrapper_80_32_inst0__I_79[31:0] = ZextWrapper_1_32_inst39__O[31:0];

  assign MuxWrapper_80_32_inst0__I_8[31:0] = ZextWrapper_2_32_inst4__O[31:0];

  assign MuxWrapper_80_32_inst0__I_9[31:0] = ZextWrapper_1_32_inst4__O[31:0];

  assign read_config_data[31:0] = MuxWrapper_80_32_inst0__O[31:0];

  assign MuxWrapper_80_32_inst0__S[0] = config_config_addr[0];

  assign MuxWrapper_80_32_inst0__S[1] = config_config_addr[1];

  assign MuxWrapper_80_32_inst0__S[2] = config_config_addr[2];

  assign MuxWrapper_80_32_inst0__S[3] = config_config_addr[3];

  assign MuxWrapper_80_32_inst0__S[4] = config_config_addr[4];

  assign MuxWrapper_80_32_inst0__S[5] = config_config_addr[5];

  assign MuxWrapper_80_32_inst0__S[6] = config_config_addr[6];

  assign reg_P_inst0__clk = clk;

  assign reg_P_inst1__clk = clk;

  assign reg_P_inst10__clk = clk;

  assign reg_P_inst11__clk = clk;

  assign reg_P_inst12__clk = clk;

  assign reg_P_inst13__clk = clk;

  assign reg_P_inst14__clk = clk;

  assign reg_P_inst15__clk = clk;

  assign reg_P_inst16__clk = clk;

  assign reg_P_inst17__clk = clk;

  assign reg_P_inst18__clk = clk;

  assign reg_P_inst19__clk = clk;

  assign reg_P_inst2__clk = clk;

  assign reg_P_inst20__clk = clk;

  assign reg_P_inst21__clk = clk;

  assign reg_P_inst22__clk = clk;

  assign reg_P_inst23__clk = clk;

  assign reg_P_inst24__clk = clk;

  assign reg_P_inst25__clk = clk;

  assign reg_P_inst26__clk = clk;

  assign reg_P_inst27__clk = clk;

  assign reg_P_inst28__clk = clk;

  assign reg_P_inst29__clk = clk;

  assign reg_P_inst3__clk = clk;

  assign reg_P_inst30__clk = clk;

  assign reg_P_inst31__clk = clk;

  assign reg_P_inst32__clk = clk;

  assign reg_P_inst33__clk = clk;

  assign reg_P_inst34__clk = clk;

  assign reg_P_inst35__clk = clk;

  assign reg_P_inst36__clk = clk;

  assign reg_P_inst37__clk = clk;

  assign reg_P_inst38__clk = clk;

  assign reg_P_inst39__clk = clk;

  assign reg_P_inst4__clk = clk;

  assign reg_P_inst5__clk = clk;

  assign reg_P_inst6__clk = clk;

  assign reg_P_inst7__clk = clk;

  assign reg_P_inst8__clk = clk;

  assign reg_P_inst9__clk = clk;


endmodule  // SB_Out_Bits_16___Out_Bits_1__

module CB_10_16_unq1 (
  input [15:0] I_0,
  input [15:0] I_1,
  input [15:0] I_2,
  input [15:0] I_3,
  input [15:0] I_4,
  input [15:0] I_5,
  input [15:0] I_6,
  input [15:0] I_7,
  input [15:0] I_8,
  input [15:0] I_9,
  output [15:0] O,
  input  clk,
  input [7:0] config_config_addr,
  input [31:0] config_config_data,
  input [0:0] config_read,
  input [0:0] config_write,
  output [31:0] read_config_data,
  input  reset
);


  wire [3:0] ConfigRegister_4_8_32_0_inst0__O;
  wire  ConfigRegister_4_8_32_0_inst0__clk;
  wire [7:0] ConfigRegister_4_8_32_0_inst0__config_addr;
  wire [31:0] ConfigRegister_4_8_32_0_inst0__config_data;
  wire  ConfigRegister_4_8_32_0_inst0__config_en;
  wire  ConfigRegister_4_8_32_0_inst0__reset;
  ConfigRegister_4_8_32_0 ConfigRegister_4_8_32_0_inst0(
    .O(ConfigRegister_4_8_32_0_inst0__O),
    .clk(ConfigRegister_4_8_32_0_inst0__clk),
    .config_addr(ConfigRegister_4_8_32_0_inst0__config_addr),
    .config_data(ConfigRegister_4_8_32_0_inst0__config_data),
    .config_en(ConfigRegister_4_8_32_0_inst0__config_en),
    .reset(ConfigRegister_4_8_32_0_inst0__reset)
  );

  wire [15:0] MuxWrapper_10_16_inst0__I_0;
  wire [15:0] MuxWrapper_10_16_inst0__I_1;
  wire [15:0] MuxWrapper_10_16_inst0__I_2;
  wire [15:0] MuxWrapper_10_16_inst0__I_3;
  wire [15:0] MuxWrapper_10_16_inst0__I_4;
  wire [15:0] MuxWrapper_10_16_inst0__I_5;
  wire [15:0] MuxWrapper_10_16_inst0__I_6;
  wire [15:0] MuxWrapper_10_16_inst0__I_7;
  wire [15:0] MuxWrapper_10_16_inst0__I_8;
  wire [15:0] MuxWrapper_10_16_inst0__I_9;
  wire [15:0] MuxWrapper_10_16_inst0__O;
  wire [3:0] MuxWrapper_10_16_inst0__S;
  MuxWrapper_10_16 MuxWrapper_10_16_inst0(
    .I_0(MuxWrapper_10_16_inst0__I_0),
    .I_1(MuxWrapper_10_16_inst0__I_1),
    .I_2(MuxWrapper_10_16_inst0__I_2),
    .I_3(MuxWrapper_10_16_inst0__I_3),
    .I_4(MuxWrapper_10_16_inst0__I_4),
    .I_5(MuxWrapper_10_16_inst0__I_5),
    .I_6(MuxWrapper_10_16_inst0__I_6),
    .I_7(MuxWrapper_10_16_inst0__I_7),
    .I_8(MuxWrapper_10_16_inst0__I_8),
    .I_9(MuxWrapper_10_16_inst0__I_9),
    .O(MuxWrapper_10_16_inst0__O),
    .S(MuxWrapper_10_16_inst0__S)
  );

  wire [3:0] ZextWrapper_4_32_inst0__I;
  wire [31:0] ZextWrapper_4_32_inst0__O;
  ZextWrapper_4_32 ZextWrapper_4_32_inst0(
    .I(ZextWrapper_4_32_inst0__I),
    .O(ZextWrapper_4_32_inst0__O)
  );

  assign MuxWrapper_10_16_inst0__S[3:0] = ConfigRegister_4_8_32_0_inst0__O[3:0];

  assign ZextWrapper_4_32_inst0__I[3:0] = ConfigRegister_4_8_32_0_inst0__O[3:0];

  assign ConfigRegister_4_8_32_0_inst0__clk = clk;

  assign ConfigRegister_4_8_32_0_inst0__config_addr[7:0] = config_config_addr[7:0];

  assign ConfigRegister_4_8_32_0_inst0__config_data[31:0] = config_config_data[31:0];

  assign ConfigRegister_4_8_32_0_inst0__config_en = config_write[0];

  assign ConfigRegister_4_8_32_0_inst0__reset = reset;

  assign MuxWrapper_10_16_inst0__I_0[15:0] = I_0[15:0];

  assign MuxWrapper_10_16_inst0__I_1[15:0] = I_1[15:0];

  assign MuxWrapper_10_16_inst0__I_2[15:0] = I_2[15:0];

  assign MuxWrapper_10_16_inst0__I_3[15:0] = I_3[15:0];

  assign MuxWrapper_10_16_inst0__I_4[15:0] = I_4[15:0];

  assign MuxWrapper_10_16_inst0__I_5[15:0] = I_5[15:0];

  assign MuxWrapper_10_16_inst0__I_6[15:0] = I_6[15:0];

  assign MuxWrapper_10_16_inst0__I_7[15:0] = I_7[15:0];

  assign MuxWrapper_10_16_inst0__I_8[15:0] = I_8[15:0];

  assign MuxWrapper_10_16_inst0__I_9[15:0] = I_9[15:0];

  assign O[15:0] = MuxWrapper_10_16_inst0__O[15:0];

  assign read_config_data[31:0] = ZextWrapper_4_32_inst0__O[31:0];


endmodule  // CB_10_16_unq1

module CB_10_16 (
  input [15:0] I_0,
  input [15:0] I_1,
  input [15:0] I_2,
  input [15:0] I_3,
  input [15:0] I_4,
  input [15:0] I_5,
  input [15:0] I_6,
  input [15:0] I_7,
  input [15:0] I_8,
  input [15:0] I_9,
  output [15:0] O,
  input  clk,
  input [7:0] config_config_addr,
  input [31:0] config_config_data,
  input [0:0] config_read,
  input [0:0] config_write,
  output [31:0] read_config_data,
  input  reset
);


  wire [3:0] ConfigRegister_4_8_32_0_inst0__O;
  wire  ConfigRegister_4_8_32_0_inst0__clk;
  wire [7:0] ConfigRegister_4_8_32_0_inst0__config_addr;
  wire [31:0] ConfigRegister_4_8_32_0_inst0__config_data;
  wire  ConfigRegister_4_8_32_0_inst0__config_en;
  wire  ConfigRegister_4_8_32_0_inst0__reset;
  ConfigRegister_4_8_32_0 ConfigRegister_4_8_32_0_inst0(
    .O(ConfigRegister_4_8_32_0_inst0__O),
    .clk(ConfigRegister_4_8_32_0_inst0__clk),
    .config_addr(ConfigRegister_4_8_32_0_inst0__config_addr),
    .config_data(ConfigRegister_4_8_32_0_inst0__config_data),
    .config_en(ConfigRegister_4_8_32_0_inst0__config_en),
    .reset(ConfigRegister_4_8_32_0_inst0__reset)
  );

  wire [15:0] MuxWrapper_10_16_inst0__I_0;
  wire [15:0] MuxWrapper_10_16_inst0__I_1;
  wire [15:0] MuxWrapper_10_16_inst0__I_2;
  wire [15:0] MuxWrapper_10_16_inst0__I_3;
  wire [15:0] MuxWrapper_10_16_inst0__I_4;
  wire [15:0] MuxWrapper_10_16_inst0__I_5;
  wire [15:0] MuxWrapper_10_16_inst0__I_6;
  wire [15:0] MuxWrapper_10_16_inst0__I_7;
  wire [15:0] MuxWrapper_10_16_inst0__I_8;
  wire [15:0] MuxWrapper_10_16_inst0__I_9;
  wire [15:0] MuxWrapper_10_16_inst0__O;
  wire [3:0] MuxWrapper_10_16_inst0__S;
  MuxWrapper_10_16 MuxWrapper_10_16_inst0(
    .I_0(MuxWrapper_10_16_inst0__I_0),
    .I_1(MuxWrapper_10_16_inst0__I_1),
    .I_2(MuxWrapper_10_16_inst0__I_2),
    .I_3(MuxWrapper_10_16_inst0__I_3),
    .I_4(MuxWrapper_10_16_inst0__I_4),
    .I_5(MuxWrapper_10_16_inst0__I_5),
    .I_6(MuxWrapper_10_16_inst0__I_6),
    .I_7(MuxWrapper_10_16_inst0__I_7),
    .I_8(MuxWrapper_10_16_inst0__I_8),
    .I_9(MuxWrapper_10_16_inst0__I_9),
    .O(MuxWrapper_10_16_inst0__O),
    .S(MuxWrapper_10_16_inst0__S)
  );

  wire [3:0] ZextWrapper_4_32_inst0__I;
  wire [31:0] ZextWrapper_4_32_inst0__O;
  ZextWrapper_4_32 ZextWrapper_4_32_inst0(
    .I(ZextWrapper_4_32_inst0__I),
    .O(ZextWrapper_4_32_inst0__O)
  );

  assign MuxWrapper_10_16_inst0__S[3:0] = ConfigRegister_4_8_32_0_inst0__O[3:0];

  assign ZextWrapper_4_32_inst0__I[3:0] = ConfigRegister_4_8_32_0_inst0__O[3:0];

  assign ConfigRegister_4_8_32_0_inst0__clk = clk;

  assign ConfigRegister_4_8_32_0_inst0__config_addr[7:0] = config_config_addr[7:0];

  assign ConfigRegister_4_8_32_0_inst0__config_data[31:0] = config_config_data[31:0];

  assign ConfigRegister_4_8_32_0_inst0__config_en = config_write[0];

  assign ConfigRegister_4_8_32_0_inst0__reset = reset;

  assign MuxWrapper_10_16_inst0__I_0[15:0] = I_0[15:0];

  assign MuxWrapper_10_16_inst0__I_1[15:0] = I_1[15:0];

  assign MuxWrapper_10_16_inst0__I_2[15:0] = I_2[15:0];

  assign MuxWrapper_10_16_inst0__I_3[15:0] = I_3[15:0];

  assign MuxWrapper_10_16_inst0__I_4[15:0] = I_4[15:0];

  assign MuxWrapper_10_16_inst0__I_5[15:0] = I_5[15:0];

  assign MuxWrapper_10_16_inst0__I_6[15:0] = I_6[15:0];

  assign MuxWrapper_10_16_inst0__I_7[15:0] = I_7[15:0];

  assign MuxWrapper_10_16_inst0__I_8[15:0] = I_8[15:0];

  assign MuxWrapper_10_16_inst0__I_9[15:0] = I_9[15:0];

  assign O[15:0] = MuxWrapper_10_16_inst0__O[15:0];

  assign read_config_data[31:0] = ZextWrapper_4_32_inst0__O[31:0];


endmodule  // CB_10_16

module CB_10_1 (
  input [0:0] I_0,
  input [0:0] I_1,
  input [0:0] I_2,
  input [0:0] I_3,
  input [0:0] I_4,
  input [0:0] I_5,
  input [0:0] I_6,
  input [0:0] I_7,
  input [0:0] I_8,
  input [0:0] I_9,
  output [0:0] O,
  input  clk,
  input [7:0] config_config_addr,
  input [31:0] config_config_data,
  input [0:0] config_read,
  input [0:0] config_write,
  output [31:0] read_config_data,
  input  reset
);


  wire [3:0] ConfigRegister_4_8_32_0_inst0__O;
  wire  ConfigRegister_4_8_32_0_inst0__clk;
  wire [7:0] ConfigRegister_4_8_32_0_inst0__config_addr;
  wire [31:0] ConfigRegister_4_8_32_0_inst0__config_data;
  wire  ConfigRegister_4_8_32_0_inst0__config_en;
  wire  ConfigRegister_4_8_32_0_inst0__reset;
  ConfigRegister_4_8_32_0 ConfigRegister_4_8_32_0_inst0(
    .O(ConfigRegister_4_8_32_0_inst0__O),
    .clk(ConfigRegister_4_8_32_0_inst0__clk),
    .config_addr(ConfigRegister_4_8_32_0_inst0__config_addr),
    .config_data(ConfigRegister_4_8_32_0_inst0__config_data),
    .config_en(ConfigRegister_4_8_32_0_inst0__config_en),
    .reset(ConfigRegister_4_8_32_0_inst0__reset)
  );

  wire [0:0] MuxWrapper_10_1_inst0__I_0;
  wire [0:0] MuxWrapper_10_1_inst0__I_1;
  wire [0:0] MuxWrapper_10_1_inst0__I_2;
  wire [0:0] MuxWrapper_10_1_inst0__I_3;
  wire [0:0] MuxWrapper_10_1_inst0__I_4;
  wire [0:0] MuxWrapper_10_1_inst0__I_5;
  wire [0:0] MuxWrapper_10_1_inst0__I_6;
  wire [0:0] MuxWrapper_10_1_inst0__I_7;
  wire [0:0] MuxWrapper_10_1_inst0__I_8;
  wire [0:0] MuxWrapper_10_1_inst0__I_9;
  wire [0:0] MuxWrapper_10_1_inst0__O;
  wire [3:0] MuxWrapper_10_1_inst0__S;
  MuxWrapper_10_1 MuxWrapper_10_1_inst0(
    .I_0(MuxWrapper_10_1_inst0__I_0),
    .I_1(MuxWrapper_10_1_inst0__I_1),
    .I_2(MuxWrapper_10_1_inst0__I_2),
    .I_3(MuxWrapper_10_1_inst0__I_3),
    .I_4(MuxWrapper_10_1_inst0__I_4),
    .I_5(MuxWrapper_10_1_inst0__I_5),
    .I_6(MuxWrapper_10_1_inst0__I_6),
    .I_7(MuxWrapper_10_1_inst0__I_7),
    .I_8(MuxWrapper_10_1_inst0__I_8),
    .I_9(MuxWrapper_10_1_inst0__I_9),
    .O(MuxWrapper_10_1_inst0__O),
    .S(MuxWrapper_10_1_inst0__S)
  );

  wire [3:0] ZextWrapper_4_32_inst0__I;
  wire [31:0] ZextWrapper_4_32_inst0__O;
  ZextWrapper_4_32 ZextWrapper_4_32_inst0(
    .I(ZextWrapper_4_32_inst0__I),
    .O(ZextWrapper_4_32_inst0__O)
  );

  assign MuxWrapper_10_1_inst0__S[3:0] = ConfigRegister_4_8_32_0_inst0__O[3:0];

  assign ZextWrapper_4_32_inst0__I[3:0] = ConfigRegister_4_8_32_0_inst0__O[3:0];

  assign ConfigRegister_4_8_32_0_inst0__clk = clk;

  assign ConfigRegister_4_8_32_0_inst0__config_addr[7:0] = config_config_addr[7:0];

  assign ConfigRegister_4_8_32_0_inst0__config_data[31:0] = config_config_data[31:0];

  assign ConfigRegister_4_8_32_0_inst0__config_en = config_write[0];

  assign ConfigRegister_4_8_32_0_inst0__reset = reset;

  assign MuxWrapper_10_1_inst0__I_0[0:0] = I_0[0:0];

  assign MuxWrapper_10_1_inst0__I_1[0:0] = I_1[0:0];

  assign MuxWrapper_10_1_inst0__I_2[0:0] = I_2[0:0];

  assign MuxWrapper_10_1_inst0__I_3[0:0] = I_3[0:0];

  assign MuxWrapper_10_1_inst0__I_4[0:0] = I_4[0:0];

  assign MuxWrapper_10_1_inst0__I_5[0:0] = I_5[0:0];

  assign MuxWrapper_10_1_inst0__I_6[0:0] = I_6[0:0];

  assign MuxWrapper_10_1_inst0__I_7[0:0] = I_7[0:0];

  assign MuxWrapper_10_1_inst0__I_8[0:0] = I_8[0:0];

  assign MuxWrapper_10_1_inst0__I_9[0:0] = I_9[0:0];

  assign O[0:0] = MuxWrapper_10_1_inst0__O[0:0];

  assign read_config_data[31:0] = ZextWrapper_4_32_inst0__O[31:0];


endmodule  // CB_10_1

module Tile_PECore (
  input  clk,
  input [31:0] config_config_addr,
  input [31:0] config_config_data,
  input [0:0] config_read,
  input [0:0] config_write,
  input [15:0] east_I_layer16_0,
  input [15:0] east_I_layer16_1,
  input [15:0] east_I_layer16_2,
  input [15:0] east_I_layer16_3,
  input [15:0] east_I_layer16_4,
  input [0:0] east_I_layer1_0,
  input [0:0] east_I_layer1_1,
  input [0:0] east_I_layer1_2,
  input [0:0] east_I_layer1_3,
  input [0:0] east_I_layer1_4,
  output [15:0] east_O_layer16_0,
  output [15:0] east_O_layer16_1,
  output [15:0] east_O_layer16_2,
  output [15:0] east_O_layer16_3,
  output [15:0] east_O_layer16_4,
  output [0:0] east_O_layer1_0,
  output [0:0] east_O_layer1_1,
  output [0:0] east_O_layer1_2,
  output [0:0] east_O_layer1_3,
  output [0:0] east_O_layer1_4,
  input [15:0] north_I_layer16_0,
  input [15:0] north_I_layer16_1,
  input [15:0] north_I_layer16_2,
  input [15:0] north_I_layer16_3,
  input [15:0] north_I_layer16_4,
  input [0:0] north_I_layer1_0,
  input [0:0] north_I_layer1_1,
  input [0:0] north_I_layer1_2,
  input [0:0] north_I_layer1_3,
  input [0:0] north_I_layer1_4,
  output [15:0] north_O_layer16_0,
  output [15:0] north_O_layer16_1,
  output [15:0] north_O_layer16_2,
  output [15:0] north_O_layer16_3,
  output [15:0] north_O_layer16_4,
  output [0:0] north_O_layer1_0,
  output [0:0] north_O_layer1_1,
  output [0:0] north_O_layer1_2,
  output [0:0] north_O_layer1_3,
  output [0:0] north_O_layer1_4,
  output [31:0] read_config_data,
  input  reset,
  input [15:0] south_I_layer16_0,
  input [15:0] south_I_layer16_1,
  input [15:0] south_I_layer16_2,
  input [15:0] south_I_layer16_3,
  input [15:0] south_I_layer16_4,
  input [0:0] south_I_layer1_0,
  input [0:0] south_I_layer1_1,
  input [0:0] south_I_layer1_2,
  input [0:0] south_I_layer1_3,
  input [0:0] south_I_layer1_4,
  output [15:0] south_O_layer16_0,
  output [15:0] south_O_layer16_1,
  output [15:0] south_O_layer16_2,
  output [15:0] south_O_layer16_3,
  output [15:0] south_O_layer16_4,
  output [0:0] south_O_layer1_0,
  output [0:0] south_O_layer1_1,
  output [0:0] south_O_layer1_2,
  output [0:0] south_O_layer1_3,
  output [0:0] south_O_layer1_4,
  input [3:0] stall,
  input [15:0] tile_id,
  input [15:0] west_I_layer16_0,
  input [15:0] west_I_layer16_1,
  input [15:0] west_I_layer16_2,
  input [15:0] west_I_layer16_3,
  input [15:0] west_I_layer16_4,
  input [0:0] west_I_layer1_0,
  input [0:0] west_I_layer1_1,
  input [0:0] west_I_layer1_2,
  input [0:0] west_I_layer1_3,
  input [0:0] west_I_layer1_4,
  output [15:0] west_O_layer16_0,
  output [15:0] west_O_layer16_1,
  output [15:0] west_O_layer16_2,
  output [15:0] west_O_layer16_3,
  output [15:0] west_O_layer16_4,
  output [0:0] west_O_layer1_0,
  output [0:0] west_O_layer1_1,
  output [0:0] west_O_layer1_2,
  output [0:0] west_O_layer1_3,
  output [0:0] west_O_layer1_4
);


  wire [15:0] CB_10_16_inst0__I_0;
  wire [15:0] CB_10_16_inst0__I_1;
  wire [15:0] CB_10_16_inst0__I_2;
  wire [15:0] CB_10_16_inst0__I_3;
  wire [15:0] CB_10_16_inst0__I_4;
  wire [15:0] CB_10_16_inst0__I_5;
  wire [15:0] CB_10_16_inst0__I_6;
  wire [15:0] CB_10_16_inst0__I_7;
  wire [15:0] CB_10_16_inst0__I_8;
  wire [15:0] CB_10_16_inst0__I_9;
  wire [15:0] CB_10_16_inst0__O;
  wire  CB_10_16_inst0__clk;
  wire [7:0] CB_10_16_inst0__config_config_addr;
  wire [31:0] CB_10_16_inst0__config_config_data;
  wire [0:0] CB_10_16_inst0__config_read;
  wire [0:0] CB_10_16_inst0__config_write;
  wire [31:0] CB_10_16_inst0__read_config_data;
  wire  CB_10_16_inst0__reset;
  CB_10_16 CB_10_16_inst0(
    .I_0(CB_10_16_inst0__I_0),
    .I_1(CB_10_16_inst0__I_1),
    .I_2(CB_10_16_inst0__I_2),
    .I_3(CB_10_16_inst0__I_3),
    .I_4(CB_10_16_inst0__I_4),
    .I_5(CB_10_16_inst0__I_5),
    .I_6(CB_10_16_inst0__I_6),
    .I_7(CB_10_16_inst0__I_7),
    .I_8(CB_10_16_inst0__I_8),
    .I_9(CB_10_16_inst0__I_9),
    .O(CB_10_16_inst0__O),
    .clk(CB_10_16_inst0__clk),
    .config_config_addr(CB_10_16_inst0__config_config_addr),
    .config_config_data(CB_10_16_inst0__config_config_data),
    .config_read(CB_10_16_inst0__config_read),
    .config_write(CB_10_16_inst0__config_write),
    .read_config_data(CB_10_16_inst0__read_config_data),
    .reset(CB_10_16_inst0__reset)
  );

  wire [15:0] CB_10_16_inst1__I_0;
  wire [15:0] CB_10_16_inst1__I_1;
  wire [15:0] CB_10_16_inst1__I_2;
  wire [15:0] CB_10_16_inst1__I_3;
  wire [15:0] CB_10_16_inst1__I_4;
  wire [15:0] CB_10_16_inst1__I_5;
  wire [15:0] CB_10_16_inst1__I_6;
  wire [15:0] CB_10_16_inst1__I_7;
  wire [15:0] CB_10_16_inst1__I_8;
  wire [15:0] CB_10_16_inst1__I_9;
  wire [15:0] CB_10_16_inst1__O;
  wire  CB_10_16_inst1__clk;
  wire [7:0] CB_10_16_inst1__config_config_addr;
  wire [31:0] CB_10_16_inst1__config_config_data;
  wire [0:0] CB_10_16_inst1__config_read;
  wire [0:0] CB_10_16_inst1__config_write;
  wire [31:0] CB_10_16_inst1__read_config_data;
  wire  CB_10_16_inst1__reset;
  CB_10_16_unq1 CB_10_16_inst1(
    .I_0(CB_10_16_inst1__I_0),
    .I_1(CB_10_16_inst1__I_1),
    .I_2(CB_10_16_inst1__I_2),
    .I_3(CB_10_16_inst1__I_3),
    .I_4(CB_10_16_inst1__I_4),
    .I_5(CB_10_16_inst1__I_5),
    .I_6(CB_10_16_inst1__I_6),
    .I_7(CB_10_16_inst1__I_7),
    .I_8(CB_10_16_inst1__I_8),
    .I_9(CB_10_16_inst1__I_9),
    .O(CB_10_16_inst1__O),
    .clk(CB_10_16_inst1__clk),
    .config_config_addr(CB_10_16_inst1__config_config_addr),
    .config_config_data(CB_10_16_inst1__config_config_data),
    .config_read(CB_10_16_inst1__config_read),
    .config_write(CB_10_16_inst1__config_write),
    .read_config_data(CB_10_16_inst1__read_config_data),
    .reset(CB_10_16_inst1__reset)
  );

  wire [0:0] CB_10_1_inst0__I_0;
  wire [0:0] CB_10_1_inst0__I_1;
  wire [0:0] CB_10_1_inst0__I_2;
  wire [0:0] CB_10_1_inst0__I_3;
  wire [0:0] CB_10_1_inst0__I_4;
  wire [0:0] CB_10_1_inst0__I_5;
  wire [0:0] CB_10_1_inst0__I_6;
  wire [0:0] CB_10_1_inst0__I_7;
  wire [0:0] CB_10_1_inst0__I_8;
  wire [0:0] CB_10_1_inst0__I_9;
  wire [0:0] CB_10_1_inst0__O;
  wire  CB_10_1_inst0__clk;
  wire [7:0] CB_10_1_inst0__config_config_addr;
  wire [31:0] CB_10_1_inst0__config_config_data;
  wire [0:0] CB_10_1_inst0__config_read;
  wire [0:0] CB_10_1_inst0__config_write;
  wire [31:0] CB_10_1_inst0__read_config_data;
  wire  CB_10_1_inst0__reset;
  CB_10_1 CB_10_1_inst0(
    .I_0(CB_10_1_inst0__I_0),
    .I_1(CB_10_1_inst0__I_1),
    .I_2(CB_10_1_inst0__I_2),
    .I_3(CB_10_1_inst0__I_3),
    .I_4(CB_10_1_inst0__I_4),
    .I_5(CB_10_1_inst0__I_5),
    .I_6(CB_10_1_inst0__I_6),
    .I_7(CB_10_1_inst0__I_7),
    .I_8(CB_10_1_inst0__I_8),
    .I_9(CB_10_1_inst0__I_9),
    .O(CB_10_1_inst0__O),
    .clk(CB_10_1_inst0__clk),
    .config_config_addr(CB_10_1_inst0__config_config_addr),
    .config_config_data(CB_10_1_inst0__config_config_data),
    .config_read(CB_10_1_inst0__config_read),
    .config_write(CB_10_1_inst0__config_write),
    .read_config_data(CB_10_1_inst0__read_config_data),
    .reset(CB_10_1_inst0__reset)
  );

  wire [0:0] CB_10_1_inst1__I_0;
  wire [0:0] CB_10_1_inst1__I_1;
  wire [0:0] CB_10_1_inst1__I_2;
  wire [0:0] CB_10_1_inst1__I_3;
  wire [0:0] CB_10_1_inst1__I_4;
  wire [0:0] CB_10_1_inst1__I_5;
  wire [0:0] CB_10_1_inst1__I_6;
  wire [0:0] CB_10_1_inst1__I_7;
  wire [0:0] CB_10_1_inst1__I_8;
  wire [0:0] CB_10_1_inst1__I_9;
  wire [0:0] CB_10_1_inst1__O;
  wire  CB_10_1_inst1__clk;
  wire [7:0] CB_10_1_inst1__config_config_addr;
  wire [31:0] CB_10_1_inst1__config_config_data;
  wire [0:0] CB_10_1_inst1__config_read;
  wire [0:0] CB_10_1_inst1__config_write;
  wire [31:0] CB_10_1_inst1__read_config_data;
  wire  CB_10_1_inst1__reset;
  CB_10_1 CB_10_1_inst1(
    .I_0(CB_10_1_inst1__I_0),
    .I_1(CB_10_1_inst1__I_1),
    .I_2(CB_10_1_inst1__I_2),
    .I_3(CB_10_1_inst1__I_3),
    .I_4(CB_10_1_inst1__I_4),
    .I_5(CB_10_1_inst1__I_5),
    .I_6(CB_10_1_inst1__I_6),
    .I_7(CB_10_1_inst1__I_7),
    .I_8(CB_10_1_inst1__I_8),
    .I_9(CB_10_1_inst1__I_9),
    .O(CB_10_1_inst1__O),
    .clk(CB_10_1_inst1__clk),
    .config_config_addr(CB_10_1_inst1__config_config_addr),
    .config_config_data(CB_10_1_inst1__config_config_data),
    .config_read(CB_10_1_inst1__config_read),
    .config_write(CB_10_1_inst1__config_write),
    .read_config_data(CB_10_1_inst1__read_config_data),
    .reset(CB_10_1_inst1__reset)
  );

  wire [0:0] CB_10_1_inst2__I_0;
  wire [0:0] CB_10_1_inst2__I_1;
  wire [0:0] CB_10_1_inst2__I_2;
  wire [0:0] CB_10_1_inst2__I_3;
  wire [0:0] CB_10_1_inst2__I_4;
  wire [0:0] CB_10_1_inst2__I_5;
  wire [0:0] CB_10_1_inst2__I_6;
  wire [0:0] CB_10_1_inst2__I_7;
  wire [0:0] CB_10_1_inst2__I_8;
  wire [0:0] CB_10_1_inst2__I_9;
  wire [0:0] CB_10_1_inst2__O;
  wire  CB_10_1_inst2__clk;
  wire [7:0] CB_10_1_inst2__config_config_addr;
  wire [31:0] CB_10_1_inst2__config_config_data;
  wire [0:0] CB_10_1_inst2__config_read;
  wire [0:0] CB_10_1_inst2__config_write;
  wire [31:0] CB_10_1_inst2__read_config_data;
  wire  CB_10_1_inst2__reset;
  CB_10_1 CB_10_1_inst2(
    .I_0(CB_10_1_inst2__I_0),
    .I_1(CB_10_1_inst2__I_1),
    .I_2(CB_10_1_inst2__I_2),
    .I_3(CB_10_1_inst2__I_3),
    .I_4(CB_10_1_inst2__I_4),
    .I_5(CB_10_1_inst2__I_5),
    .I_6(CB_10_1_inst2__I_6),
    .I_7(CB_10_1_inst2__I_7),
    .I_8(CB_10_1_inst2__I_8),
    .I_9(CB_10_1_inst2__I_9),
    .O(CB_10_1_inst2__O),
    .clk(CB_10_1_inst2__clk),
    .config_config_addr(CB_10_1_inst2__config_config_addr),
    .config_config_data(CB_10_1_inst2__config_config_data),
    .config_read(CB_10_1_inst2__config_read),
    .config_write(CB_10_1_inst2__config_write),
    .read_config_data(CB_10_1_inst2__read_config_data),
    .reset(CB_10_1_inst2__reset)
  );

  wire [7:0] Decode08_inst0__I;
  wire  Decode08_inst0__O;
  Decode08 Decode08_inst0(
    .I(Decode08_inst0__I),
    .O(Decode08_inst0__O)
  );

  wire [7:0] Decode18_inst0__I;
  wire  Decode18_inst0__O;
  Decode18 Decode18_inst0(
    .I(Decode18_inst0__I),
    .O(Decode18_inst0__O)
  );

  wire [7:0] Decode28_inst0__I;
  wire  Decode28_inst0__O;
  Decode28 Decode28_inst0(
    .I(Decode28_inst0__I),
    .O(Decode28_inst0__O)
  );

  wire [7:0] Decode38_inst0__I;
  wire  Decode38_inst0__O;
  Decode38 Decode38_inst0(
    .I(Decode38_inst0__I),
    .O(Decode38_inst0__O)
  );

  wire [7:0] Decode48_inst0__I;
  wire  Decode48_inst0__O;
  Decode48 Decode48_inst0(
    .I(Decode48_inst0__I),
    .O(Decode48_inst0__O)
  );

  wire [7:0] Decode58_inst0__I;
  wire  Decode58_inst0__O;
  Decode58 Decode58_inst0(
    .I(Decode58_inst0__I),
    .O(Decode58_inst0__O)
  );

  wire [7:0] Decode68_inst0__I;
  wire  Decode68_inst0__O;
  Decode68 Decode68_inst0(
    .I(Decode68_inst0__I),
    .O(Decode68_inst0__O)
  );

  wire [0:0] MuxWithDefaultWrapper_7_32_8_0_inst0__EN;
  wire [31:0] MuxWithDefaultWrapper_7_32_8_0_inst0__I_0;
  wire [31:0] MuxWithDefaultWrapper_7_32_8_0_inst0__I_1;
  wire [31:0] MuxWithDefaultWrapper_7_32_8_0_inst0__I_2;
  wire [31:0] MuxWithDefaultWrapper_7_32_8_0_inst0__I_3;
  wire [31:0] MuxWithDefaultWrapper_7_32_8_0_inst0__I_4;
  wire [31:0] MuxWithDefaultWrapper_7_32_8_0_inst0__I_5;
  wire [31:0] MuxWithDefaultWrapper_7_32_8_0_inst0__I_6;
  wire [31:0] MuxWithDefaultWrapper_7_32_8_0_inst0__O;
  wire [7:0] MuxWithDefaultWrapper_7_32_8_0_inst0__S;
  MuxWithDefaultWrapper_7_32_8_0 MuxWithDefaultWrapper_7_32_8_0_inst0(
    .EN(MuxWithDefaultWrapper_7_32_8_0_inst0__EN),
    .I_0(MuxWithDefaultWrapper_7_32_8_0_inst0__I_0),
    .I_1(MuxWithDefaultWrapper_7_32_8_0_inst0__I_1),
    .I_2(MuxWithDefaultWrapper_7_32_8_0_inst0__I_2),
    .I_3(MuxWithDefaultWrapper_7_32_8_0_inst0__I_3),
    .I_4(MuxWithDefaultWrapper_7_32_8_0_inst0__I_4),
    .I_5(MuxWithDefaultWrapper_7_32_8_0_inst0__I_5),
    .I_6(MuxWithDefaultWrapper_7_32_8_0_inst0__I_6),
    .O(MuxWithDefaultWrapper_7_32_8_0_inst0__O),
    .S(MuxWithDefaultWrapper_7_32_8_0_inst0__S)
  );

  wire [0:0] PECore_inst0__bit0;
  wire [0:0] PECore_inst0__bit1;
  wire [0:0] PECore_inst0__bit2;
  wire  PECore_inst0__clk;
  wire [7:0] PECore_inst0__config_config_addr;
  wire [31:0] PECore_inst0__config_config_data;
  wire [0:0] PECore_inst0__config_read;
  wire [0:0] PECore_inst0__config_write;
  wire [15:0] PECore_inst0__data0;
  wire [15:0] PECore_inst0__data1;
  wire [31:0] PECore_inst0__read_config_data;
  wire [15:0] PECore_inst0__res;
  wire [0:0] PECore_inst0__res_p;
  wire  PECore_inst0__reset;
  wire [3:0] PECore_inst0__stall;
  PECore PECore_inst0(
    .bit0(PECore_inst0__bit0),
    .bit1(PECore_inst0__bit1),
    .bit2(PECore_inst0__bit2),
    .clk(PECore_inst0__clk),
    .config_config_addr(PECore_inst0__config_config_addr),
    .config_config_data(PECore_inst0__config_config_data),
    .config_read(PECore_inst0__config_read),
    .config_write(PECore_inst0__config_write),
    .data0(PECore_inst0__data0),
    .data1(PECore_inst0__data1),
    .read_config_data(PECore_inst0__read_config_data),
    .res(PECore_inst0__res),
    .res_p(PECore_inst0__res_p),
    .reset(PECore_inst0__reset),
    .stall(PECore_inst0__stall)
  );

  wire  SB_Out_Bits_16___Out_Bits_1___inst0__clk;
  wire [7:0] SB_Out_Bits_16___Out_Bits_1___inst0__config_config_addr;
  wire [31:0] SB_Out_Bits_16___Out_Bits_1___inst0__config_config_data;
  wire [0:0] SB_Out_Bits_16___Out_Bits_1___inst0__config_read;
  wire [0:0] SB_Out_Bits_16___Out_Bits_1___inst0__config_write;
  wire [15:0] SB_Out_Bits_16___Out_Bits_1___inst0__east_I_layer16_0;
  wire [15:0] SB_Out_Bits_16___Out_Bits_1___inst0__east_I_layer16_1;
  wire [15:0] SB_Out_Bits_16___Out_Bits_1___inst0__east_I_layer16_2;
  wire [15:0] SB_Out_Bits_16___Out_Bits_1___inst0__east_I_layer16_3;
  wire [15:0] SB_Out_Bits_16___Out_Bits_1___inst0__east_I_layer16_4;
  wire [0:0] SB_Out_Bits_16___Out_Bits_1___inst0__east_I_layer1_0;
  wire [0:0] SB_Out_Bits_16___Out_Bits_1___inst0__east_I_layer1_1;
  wire [0:0] SB_Out_Bits_16___Out_Bits_1___inst0__east_I_layer1_2;
  wire [0:0] SB_Out_Bits_16___Out_Bits_1___inst0__east_I_layer1_3;
  wire [0:0] SB_Out_Bits_16___Out_Bits_1___inst0__east_I_layer1_4;
  wire [15:0] SB_Out_Bits_16___Out_Bits_1___inst0__east_O_layer16_0;
  wire [15:0] SB_Out_Bits_16___Out_Bits_1___inst0__east_O_layer16_1;
  wire [15:0] SB_Out_Bits_16___Out_Bits_1___inst0__east_O_layer16_2;
  wire [15:0] SB_Out_Bits_16___Out_Bits_1___inst0__east_O_layer16_3;
  wire [15:0] SB_Out_Bits_16___Out_Bits_1___inst0__east_O_layer16_4;
  wire [0:0] SB_Out_Bits_16___Out_Bits_1___inst0__east_O_layer1_0;
  wire [0:0] SB_Out_Bits_16___Out_Bits_1___inst0__east_O_layer1_1;
  wire [0:0] SB_Out_Bits_16___Out_Bits_1___inst0__east_O_layer1_2;
  wire [0:0] SB_Out_Bits_16___Out_Bits_1___inst0__east_O_layer1_3;
  wire [0:0] SB_Out_Bits_16___Out_Bits_1___inst0__east_O_layer1_4;
  wire [15:0] SB_Out_Bits_16___Out_Bits_1___inst0__north_I_layer16_0;
  wire [15:0] SB_Out_Bits_16___Out_Bits_1___inst0__north_I_layer16_1;
  wire [15:0] SB_Out_Bits_16___Out_Bits_1___inst0__north_I_layer16_2;
  wire [15:0] SB_Out_Bits_16___Out_Bits_1___inst0__north_I_layer16_3;
  wire [15:0] SB_Out_Bits_16___Out_Bits_1___inst0__north_I_layer16_4;
  wire [0:0] SB_Out_Bits_16___Out_Bits_1___inst0__north_I_layer1_0;
  wire [0:0] SB_Out_Bits_16___Out_Bits_1___inst0__north_I_layer1_1;
  wire [0:0] SB_Out_Bits_16___Out_Bits_1___inst0__north_I_layer1_2;
  wire [0:0] SB_Out_Bits_16___Out_Bits_1___inst0__north_I_layer1_3;
  wire [0:0] SB_Out_Bits_16___Out_Bits_1___inst0__north_I_layer1_4;
  wire [15:0] SB_Out_Bits_16___Out_Bits_1___inst0__north_O_layer16_0;
  wire [15:0] SB_Out_Bits_16___Out_Bits_1___inst0__north_O_layer16_1;
  wire [15:0] SB_Out_Bits_16___Out_Bits_1___inst0__north_O_layer16_2;
  wire [15:0] SB_Out_Bits_16___Out_Bits_1___inst0__north_O_layer16_3;
  wire [15:0] SB_Out_Bits_16___Out_Bits_1___inst0__north_O_layer16_4;
  wire [0:0] SB_Out_Bits_16___Out_Bits_1___inst0__north_O_layer1_0;
  wire [0:0] SB_Out_Bits_16___Out_Bits_1___inst0__north_O_layer1_1;
  wire [0:0] SB_Out_Bits_16___Out_Bits_1___inst0__north_O_layer1_2;
  wire [0:0] SB_Out_Bits_16___Out_Bits_1___inst0__north_O_layer1_3;
  wire [0:0] SB_Out_Bits_16___Out_Bits_1___inst0__north_O_layer1_4;
  wire [31:0] SB_Out_Bits_16___Out_Bits_1___inst0__read_config_data;
  wire [15:0] SB_Out_Bits_16___Out_Bits_1___inst0__res;
  wire [0:0] SB_Out_Bits_16___Out_Bits_1___inst0__res_p;
  wire  SB_Out_Bits_16___Out_Bits_1___inst0__reset;
  wire [15:0] SB_Out_Bits_16___Out_Bits_1___inst0__south_I_layer16_0;
  wire [15:0] SB_Out_Bits_16___Out_Bits_1___inst0__south_I_layer16_1;
  wire [15:0] SB_Out_Bits_16___Out_Bits_1___inst0__south_I_layer16_2;
  wire [15:0] SB_Out_Bits_16___Out_Bits_1___inst0__south_I_layer16_3;
  wire [15:0] SB_Out_Bits_16___Out_Bits_1___inst0__south_I_layer16_4;
  wire [0:0] SB_Out_Bits_16___Out_Bits_1___inst0__south_I_layer1_0;
  wire [0:0] SB_Out_Bits_16___Out_Bits_1___inst0__south_I_layer1_1;
  wire [0:0] SB_Out_Bits_16___Out_Bits_1___inst0__south_I_layer1_2;
  wire [0:0] SB_Out_Bits_16___Out_Bits_1___inst0__south_I_layer1_3;
  wire [0:0] SB_Out_Bits_16___Out_Bits_1___inst0__south_I_layer1_4;
  wire [15:0] SB_Out_Bits_16___Out_Bits_1___inst0__south_O_layer16_0;
  wire [15:0] SB_Out_Bits_16___Out_Bits_1___inst0__south_O_layer16_1;
  wire [15:0] SB_Out_Bits_16___Out_Bits_1___inst0__south_O_layer16_2;
  wire [15:0] SB_Out_Bits_16___Out_Bits_1___inst0__south_O_layer16_3;
  wire [15:0] SB_Out_Bits_16___Out_Bits_1___inst0__south_O_layer16_4;
  wire [0:0] SB_Out_Bits_16___Out_Bits_1___inst0__south_O_layer1_0;
  wire [0:0] SB_Out_Bits_16___Out_Bits_1___inst0__south_O_layer1_1;
  wire [0:0] SB_Out_Bits_16___Out_Bits_1___inst0__south_O_layer1_2;
  wire [0:0] SB_Out_Bits_16___Out_Bits_1___inst0__south_O_layer1_3;
  wire [0:0] SB_Out_Bits_16___Out_Bits_1___inst0__south_O_layer1_4;
  wire [15:0] SB_Out_Bits_16___Out_Bits_1___inst0__west_I_layer16_0;
  wire [15:0] SB_Out_Bits_16___Out_Bits_1___inst0__west_I_layer16_1;
  wire [15:0] SB_Out_Bits_16___Out_Bits_1___inst0__west_I_layer16_2;
  wire [15:0] SB_Out_Bits_16___Out_Bits_1___inst0__west_I_layer16_3;
  wire [15:0] SB_Out_Bits_16___Out_Bits_1___inst0__west_I_layer16_4;
  wire [0:0] SB_Out_Bits_16___Out_Bits_1___inst0__west_I_layer1_0;
  wire [0:0] SB_Out_Bits_16___Out_Bits_1___inst0__west_I_layer1_1;
  wire [0:0] SB_Out_Bits_16___Out_Bits_1___inst0__west_I_layer1_2;
  wire [0:0] SB_Out_Bits_16___Out_Bits_1___inst0__west_I_layer1_3;
  wire [0:0] SB_Out_Bits_16___Out_Bits_1___inst0__west_I_layer1_4;
  wire [15:0] SB_Out_Bits_16___Out_Bits_1___inst0__west_O_layer16_0;
  wire [15:0] SB_Out_Bits_16___Out_Bits_1___inst0__west_O_layer16_1;
  wire [15:0] SB_Out_Bits_16___Out_Bits_1___inst0__west_O_layer16_2;
  wire [15:0] SB_Out_Bits_16___Out_Bits_1___inst0__west_O_layer16_3;
  wire [15:0] SB_Out_Bits_16___Out_Bits_1___inst0__west_O_layer16_4;
  wire [0:0] SB_Out_Bits_16___Out_Bits_1___inst0__west_O_layer1_0;
  wire [0:0] SB_Out_Bits_16___Out_Bits_1___inst0__west_O_layer1_1;
  wire [0:0] SB_Out_Bits_16___Out_Bits_1___inst0__west_O_layer1_2;
  wire [0:0] SB_Out_Bits_16___Out_Bits_1___inst0__west_O_layer1_3;
  wire [0:0] SB_Out_Bits_16___Out_Bits_1___inst0__west_O_layer1_4;
  SB_Out_Bits_16___Out_Bits_1__ SB_Out_Bits_16___Out_Bits_1___inst0(
    .clk(SB_Out_Bits_16___Out_Bits_1___inst0__clk),
    .config_config_addr(SB_Out_Bits_16___Out_Bits_1___inst0__config_config_addr),
    .config_config_data(SB_Out_Bits_16___Out_Bits_1___inst0__config_config_data),
    .config_read(SB_Out_Bits_16___Out_Bits_1___inst0__config_read),
    .config_write(SB_Out_Bits_16___Out_Bits_1___inst0__config_write),
    .east_I_layer16_0(SB_Out_Bits_16___Out_Bits_1___inst0__east_I_layer16_0),
    .east_I_layer16_1(SB_Out_Bits_16___Out_Bits_1___inst0__east_I_layer16_1),
    .east_I_layer16_2(SB_Out_Bits_16___Out_Bits_1___inst0__east_I_layer16_2),
    .east_I_layer16_3(SB_Out_Bits_16___Out_Bits_1___inst0__east_I_layer16_3),
    .east_I_layer16_4(SB_Out_Bits_16___Out_Bits_1___inst0__east_I_layer16_4),
    .east_I_layer1_0(SB_Out_Bits_16___Out_Bits_1___inst0__east_I_layer1_0),
    .east_I_layer1_1(SB_Out_Bits_16___Out_Bits_1___inst0__east_I_layer1_1),
    .east_I_layer1_2(SB_Out_Bits_16___Out_Bits_1___inst0__east_I_layer1_2),
    .east_I_layer1_3(SB_Out_Bits_16___Out_Bits_1___inst0__east_I_layer1_3),
    .east_I_layer1_4(SB_Out_Bits_16___Out_Bits_1___inst0__east_I_layer1_4),
    .east_O_layer16_0(SB_Out_Bits_16___Out_Bits_1___inst0__east_O_layer16_0),
    .east_O_layer16_1(SB_Out_Bits_16___Out_Bits_1___inst0__east_O_layer16_1),
    .east_O_layer16_2(SB_Out_Bits_16___Out_Bits_1___inst0__east_O_layer16_2),
    .east_O_layer16_3(SB_Out_Bits_16___Out_Bits_1___inst0__east_O_layer16_3),
    .east_O_layer16_4(SB_Out_Bits_16___Out_Bits_1___inst0__east_O_layer16_4),
    .east_O_layer1_0(SB_Out_Bits_16___Out_Bits_1___inst0__east_O_layer1_0),
    .east_O_layer1_1(SB_Out_Bits_16___Out_Bits_1___inst0__east_O_layer1_1),
    .east_O_layer1_2(SB_Out_Bits_16___Out_Bits_1___inst0__east_O_layer1_2),
    .east_O_layer1_3(SB_Out_Bits_16___Out_Bits_1___inst0__east_O_layer1_3),
    .east_O_layer1_4(SB_Out_Bits_16___Out_Bits_1___inst0__east_O_layer1_4),
    .north_I_layer16_0(SB_Out_Bits_16___Out_Bits_1___inst0__north_I_layer16_0),
    .north_I_layer16_1(SB_Out_Bits_16___Out_Bits_1___inst0__north_I_layer16_1),
    .north_I_layer16_2(SB_Out_Bits_16___Out_Bits_1___inst0__north_I_layer16_2),
    .north_I_layer16_3(SB_Out_Bits_16___Out_Bits_1___inst0__north_I_layer16_3),
    .north_I_layer16_4(SB_Out_Bits_16___Out_Bits_1___inst0__north_I_layer16_4),
    .north_I_layer1_0(SB_Out_Bits_16___Out_Bits_1___inst0__north_I_layer1_0),
    .north_I_layer1_1(SB_Out_Bits_16___Out_Bits_1___inst0__north_I_layer1_1),
    .north_I_layer1_2(SB_Out_Bits_16___Out_Bits_1___inst0__north_I_layer1_2),
    .north_I_layer1_3(SB_Out_Bits_16___Out_Bits_1___inst0__north_I_layer1_3),
    .north_I_layer1_4(SB_Out_Bits_16___Out_Bits_1___inst0__north_I_layer1_4),
    .north_O_layer16_0(SB_Out_Bits_16___Out_Bits_1___inst0__north_O_layer16_0),
    .north_O_layer16_1(SB_Out_Bits_16___Out_Bits_1___inst0__north_O_layer16_1),
    .north_O_layer16_2(SB_Out_Bits_16___Out_Bits_1___inst0__north_O_layer16_2),
    .north_O_layer16_3(SB_Out_Bits_16___Out_Bits_1___inst0__north_O_layer16_3),
    .north_O_layer16_4(SB_Out_Bits_16___Out_Bits_1___inst0__north_O_layer16_4),
    .north_O_layer1_0(SB_Out_Bits_16___Out_Bits_1___inst0__north_O_layer1_0),
    .north_O_layer1_1(SB_Out_Bits_16___Out_Bits_1___inst0__north_O_layer1_1),
    .north_O_layer1_2(SB_Out_Bits_16___Out_Bits_1___inst0__north_O_layer1_2),
    .north_O_layer1_3(SB_Out_Bits_16___Out_Bits_1___inst0__north_O_layer1_3),
    .north_O_layer1_4(SB_Out_Bits_16___Out_Bits_1___inst0__north_O_layer1_4),
    .read_config_data(SB_Out_Bits_16___Out_Bits_1___inst0__read_config_data),
    .res(SB_Out_Bits_16___Out_Bits_1___inst0__res),
    .res_p(SB_Out_Bits_16___Out_Bits_1___inst0__res_p),
    .reset(SB_Out_Bits_16___Out_Bits_1___inst0__reset),
    .south_I_layer16_0(SB_Out_Bits_16___Out_Bits_1___inst0__south_I_layer16_0),
    .south_I_layer16_1(SB_Out_Bits_16___Out_Bits_1___inst0__south_I_layer16_1),
    .south_I_layer16_2(SB_Out_Bits_16___Out_Bits_1___inst0__south_I_layer16_2),
    .south_I_layer16_3(SB_Out_Bits_16___Out_Bits_1___inst0__south_I_layer16_3),
    .south_I_layer16_4(SB_Out_Bits_16___Out_Bits_1___inst0__south_I_layer16_4),
    .south_I_layer1_0(SB_Out_Bits_16___Out_Bits_1___inst0__south_I_layer1_0),
    .south_I_layer1_1(SB_Out_Bits_16___Out_Bits_1___inst0__south_I_layer1_1),
    .south_I_layer1_2(SB_Out_Bits_16___Out_Bits_1___inst0__south_I_layer1_2),
    .south_I_layer1_3(SB_Out_Bits_16___Out_Bits_1___inst0__south_I_layer1_3),
    .south_I_layer1_4(SB_Out_Bits_16___Out_Bits_1___inst0__south_I_layer1_4),
    .south_O_layer16_0(SB_Out_Bits_16___Out_Bits_1___inst0__south_O_layer16_0),
    .south_O_layer16_1(SB_Out_Bits_16___Out_Bits_1___inst0__south_O_layer16_1),
    .south_O_layer16_2(SB_Out_Bits_16___Out_Bits_1___inst0__south_O_layer16_2),
    .south_O_layer16_3(SB_Out_Bits_16___Out_Bits_1___inst0__south_O_layer16_3),
    .south_O_layer16_4(SB_Out_Bits_16___Out_Bits_1___inst0__south_O_layer16_4),
    .south_O_layer1_0(SB_Out_Bits_16___Out_Bits_1___inst0__south_O_layer1_0),
    .south_O_layer1_1(SB_Out_Bits_16___Out_Bits_1___inst0__south_O_layer1_1),
    .south_O_layer1_2(SB_Out_Bits_16___Out_Bits_1___inst0__south_O_layer1_2),
    .south_O_layer1_3(SB_Out_Bits_16___Out_Bits_1___inst0__south_O_layer1_3),
    .south_O_layer1_4(SB_Out_Bits_16___Out_Bits_1___inst0__south_O_layer1_4),
    .west_I_layer16_0(SB_Out_Bits_16___Out_Bits_1___inst0__west_I_layer16_0),
    .west_I_layer16_1(SB_Out_Bits_16___Out_Bits_1___inst0__west_I_layer16_1),
    .west_I_layer16_2(SB_Out_Bits_16___Out_Bits_1___inst0__west_I_layer16_2),
    .west_I_layer16_3(SB_Out_Bits_16___Out_Bits_1___inst0__west_I_layer16_3),
    .west_I_layer16_4(SB_Out_Bits_16___Out_Bits_1___inst0__west_I_layer16_4),
    .west_I_layer1_0(SB_Out_Bits_16___Out_Bits_1___inst0__west_I_layer1_0),
    .west_I_layer1_1(SB_Out_Bits_16___Out_Bits_1___inst0__west_I_layer1_1),
    .west_I_layer1_2(SB_Out_Bits_16___Out_Bits_1___inst0__west_I_layer1_2),
    .west_I_layer1_3(SB_Out_Bits_16___Out_Bits_1___inst0__west_I_layer1_3),
    .west_I_layer1_4(SB_Out_Bits_16___Out_Bits_1___inst0__west_I_layer1_4),
    .west_O_layer16_0(SB_Out_Bits_16___Out_Bits_1___inst0__west_O_layer16_0),
    .west_O_layer16_1(SB_Out_Bits_16___Out_Bits_1___inst0__west_O_layer16_1),
    .west_O_layer16_2(SB_Out_Bits_16___Out_Bits_1___inst0__west_O_layer16_2),
    .west_O_layer16_3(SB_Out_Bits_16___Out_Bits_1___inst0__west_O_layer16_3),
    .west_O_layer16_4(SB_Out_Bits_16___Out_Bits_1___inst0__west_O_layer16_4),
    .west_O_layer1_0(SB_Out_Bits_16___Out_Bits_1___inst0__west_O_layer1_0),
    .west_O_layer1_1(SB_Out_Bits_16___Out_Bits_1___inst0__west_O_layer1_1),
    .west_O_layer1_2(SB_Out_Bits_16___Out_Bits_1___inst0__west_O_layer1_2),
    .west_O_layer1_3(SB_Out_Bits_16___Out_Bits_1___inst0__west_O_layer1_3),
    .west_O_layer1_4(SB_Out_Bits_16___Out_Bits_1___inst0__west_O_layer1_4)
  );

  wire  and_inst0__in0;
  wire  and_inst0__in1;
  wire  and_inst0__out;
  corebit_and and_inst0(
    .in0(and_inst0__in0),
    .in1(and_inst0__in1),
    .out(and_inst0__out)
  );

  wire  and_inst1__in0;
  wire  and_inst1__in1;
  wire  and_inst1__out;
  corebit_and and_inst1(
    .in0(and_inst1__in0),
    .in1(and_inst1__in1),
    .out(and_inst1__out)
  );

  wire  and_inst2__in0;
  wire  and_inst2__in1;
  wire  and_inst2__out;
  corebit_and and_inst2(
    .in0(and_inst2__in0),
    .in1(and_inst2__in1),
    .out(and_inst2__out)
  );

  wire  and_inst3__in0;
  wire  and_inst3__in1;
  wire  and_inst3__out;
  corebit_and and_inst3(
    .in0(and_inst3__in0),
    .in1(and_inst3__in1),
    .out(and_inst3__out)
  );

  wire  and_inst4__in0;
  wire  and_inst4__in1;
  wire  and_inst4__out;
  corebit_and and_inst4(
    .in0(and_inst4__in0),
    .in1(and_inst4__in1),
    .out(and_inst4__out)
  );

  wire  and_inst5__in0;
  wire  and_inst5__in1;
  wire  and_inst5__out;
  corebit_and and_inst5(
    .in0(and_inst5__in0),
    .in1(and_inst5__in1),
    .out(and_inst5__out)
  );

  wire  and_inst6__in0;
  wire  and_inst6__in1;
  wire  and_inst6__out;
  corebit_and and_inst6(
    .in0(and_inst6__in0),
    .in1(and_inst6__in1),
    .out(and_inst6__out)
  );

  wire  and_inst7__in0;
  wire  and_inst7__in1;
  wire  and_inst7__out;
  corebit_and and_inst7(
    .in0(and_inst7__in0),
    .in1(and_inst7__in1),
    .out(and_inst7__out)
  );

  wire  and_inst8__in0;
  wire  and_inst8__in1;
  wire  and_inst8__out;
  corebit_and and_inst8(
    .in0(and_inst8__in0),
    .in1(and_inst8__in1),
    .out(and_inst8__out)
  );

  // Instancing generated Module: coreir.eq(width:16)
  wire [15:0] coreir_eq_16_inst0__in0;
  wire [15:0] coreir_eq_16_inst0__in1;
  wire  coreir_eq_16_inst0__out;
  coreir_eq #(.width(16)) coreir_eq_16_inst0(
    .in0(coreir_eq_16_inst0__in0),
    .in1(coreir_eq_16_inst0__in1),
    .out(coreir_eq_16_inst0__out)
  );

  assign CB_10_16_inst0__I_0[15:0] = north_I_layer16_0[15:0];

  assign CB_10_16_inst0__I_1[15:0] = north_I_layer16_1[15:0];

  assign CB_10_16_inst0__I_2[15:0] = north_I_layer16_2[15:0];

  assign CB_10_16_inst0__I_3[15:0] = north_I_layer16_3[15:0];

  assign CB_10_16_inst0__I_4[15:0] = north_I_layer16_4[15:0];

  assign CB_10_16_inst0__I_5[15:0] = SB_Out_Bits_16___Out_Bits_1___inst0__north_O_layer16_0[15:0];

  assign CB_10_16_inst0__I_6[15:0] = SB_Out_Bits_16___Out_Bits_1___inst0__north_O_layer16_1[15:0];

  assign CB_10_16_inst0__I_7[15:0] = SB_Out_Bits_16___Out_Bits_1___inst0__north_O_layer16_2[15:0];

  assign CB_10_16_inst0__I_8[15:0] = SB_Out_Bits_16___Out_Bits_1___inst0__north_O_layer16_3[15:0];

  assign CB_10_16_inst0__I_9[15:0] = SB_Out_Bits_16___Out_Bits_1___inst0__north_O_layer16_4[15:0];

  assign PECore_inst0__data0[15:0] = CB_10_16_inst0__O[15:0];

  assign CB_10_16_inst0__clk = clk;

  assign CB_10_16_inst0__config_config_addr[0] = config_config_addr[24];

  assign CB_10_16_inst0__config_config_addr[1] = config_config_addr[25];

  assign CB_10_16_inst0__config_config_addr[2] = config_config_addr[26];

  assign CB_10_16_inst0__config_config_addr[3] = config_config_addr[27];

  assign CB_10_16_inst0__config_config_addr[4] = config_config_addr[28];

  assign CB_10_16_inst0__config_config_addr[5] = config_config_addr[29];

  assign CB_10_16_inst0__config_config_addr[6] = config_config_addr[30];

  assign CB_10_16_inst0__config_config_addr[7] = config_config_addr[31];

  assign CB_10_16_inst0__config_config_data[31:0] = config_config_data[31:0];

  assign CB_10_16_inst0__config_read[0:0] = config_read[0:0];

  assign CB_10_16_inst0__config_write[0] = and_inst4__out;

  assign MuxWithDefaultWrapper_7_32_8_0_inst0__I_2[31:0] = CB_10_16_inst0__read_config_data[31:0];

  assign CB_10_16_inst0__reset = reset;

  assign CB_10_16_inst1__I_0[15:0] = west_I_layer16_0[15:0];

  assign CB_10_16_inst1__I_1[15:0] = west_I_layer16_1[15:0];

  assign CB_10_16_inst1__I_2[15:0] = west_I_layer16_2[15:0];

  assign CB_10_16_inst1__I_3[15:0] = west_I_layer16_3[15:0];

  assign CB_10_16_inst1__I_4[15:0] = west_I_layer16_4[15:0];

  assign CB_10_16_inst1__I_5[15:0] = SB_Out_Bits_16___Out_Bits_1___inst0__west_O_layer16_0[15:0];

  assign CB_10_16_inst1__I_6[15:0] = SB_Out_Bits_16___Out_Bits_1___inst0__west_O_layer16_1[15:0];

  assign CB_10_16_inst1__I_7[15:0] = SB_Out_Bits_16___Out_Bits_1___inst0__west_O_layer16_2[15:0];

  assign CB_10_16_inst1__I_8[15:0] = SB_Out_Bits_16___Out_Bits_1___inst0__west_O_layer16_3[15:0];

  assign CB_10_16_inst1__I_9[15:0] = SB_Out_Bits_16___Out_Bits_1___inst0__west_O_layer16_4[15:0];

  assign PECore_inst0__data1[15:0] = CB_10_16_inst1__O[15:0];

  assign CB_10_16_inst1__clk = clk;

  assign CB_10_16_inst1__config_config_addr[0] = config_config_addr[24];

  assign CB_10_16_inst1__config_config_addr[1] = config_config_addr[25];

  assign CB_10_16_inst1__config_config_addr[2] = config_config_addr[26];

  assign CB_10_16_inst1__config_config_addr[3] = config_config_addr[27];

  assign CB_10_16_inst1__config_config_addr[4] = config_config_addr[28];

  assign CB_10_16_inst1__config_config_addr[5] = config_config_addr[29];

  assign CB_10_16_inst1__config_config_addr[6] = config_config_addr[30];

  assign CB_10_16_inst1__config_config_addr[7] = config_config_addr[31];

  assign CB_10_16_inst1__config_config_data[31:0] = config_config_data[31:0];

  assign CB_10_16_inst1__config_read[0:0] = config_read[0:0];

  assign CB_10_16_inst1__config_write[0] = and_inst5__out;

  assign MuxWithDefaultWrapper_7_32_8_0_inst0__I_3[31:0] = CB_10_16_inst1__read_config_data[31:0];

  assign CB_10_16_inst1__reset = reset;

  assign CB_10_1_inst0__I_0[0:0] = north_I_layer1_0[0:0];

  assign CB_10_1_inst0__I_1[0:0] = north_I_layer1_1[0:0];

  assign CB_10_1_inst0__I_2[0:0] = north_I_layer1_2[0:0];

  assign CB_10_1_inst0__I_3[0:0] = north_I_layer1_3[0:0];

  assign CB_10_1_inst0__I_4[0:0] = north_I_layer1_4[0:0];

  assign CB_10_1_inst0__I_5[0:0] = SB_Out_Bits_16___Out_Bits_1___inst0__north_O_layer1_0[0:0];

  assign CB_10_1_inst0__I_6[0:0] = SB_Out_Bits_16___Out_Bits_1___inst0__north_O_layer1_1[0:0];

  assign CB_10_1_inst0__I_7[0:0] = SB_Out_Bits_16___Out_Bits_1___inst0__north_O_layer1_2[0:0];

  assign CB_10_1_inst0__I_8[0:0] = SB_Out_Bits_16___Out_Bits_1___inst0__north_O_layer1_3[0:0];

  assign CB_10_1_inst0__I_9[0:0] = SB_Out_Bits_16___Out_Bits_1___inst0__north_O_layer1_4[0:0];

  assign PECore_inst0__bit0[0:0] = CB_10_1_inst0__O[0:0];

  assign CB_10_1_inst0__clk = clk;

  assign CB_10_1_inst0__config_config_addr[0] = config_config_addr[24];

  assign CB_10_1_inst0__config_config_addr[1] = config_config_addr[25];

  assign CB_10_1_inst0__config_config_addr[2] = config_config_addr[26];

  assign CB_10_1_inst0__config_config_addr[3] = config_config_addr[27];

  assign CB_10_1_inst0__config_config_addr[4] = config_config_addr[28];

  assign CB_10_1_inst0__config_config_addr[5] = config_config_addr[29];

  assign CB_10_1_inst0__config_config_addr[6] = config_config_addr[30];

  assign CB_10_1_inst0__config_config_addr[7] = config_config_addr[31];

  assign CB_10_1_inst0__config_config_data[31:0] = config_config_data[31:0];

  assign CB_10_1_inst0__config_read[0:0] = config_read[0:0];

  assign CB_10_1_inst0__config_write[0] = and_inst6__out;

  assign MuxWithDefaultWrapper_7_32_8_0_inst0__I_4[31:0] = CB_10_1_inst0__read_config_data[31:0];

  assign CB_10_1_inst0__reset = reset;

  assign CB_10_1_inst1__I_0[0:0] = west_I_layer1_0[0:0];

  assign CB_10_1_inst1__I_1[0:0] = west_I_layer1_1[0:0];

  assign CB_10_1_inst1__I_2[0:0] = west_I_layer1_2[0:0];

  assign CB_10_1_inst1__I_3[0:0] = west_I_layer1_3[0:0];

  assign CB_10_1_inst1__I_4[0:0] = west_I_layer1_4[0:0];

  assign CB_10_1_inst1__I_5[0:0] = SB_Out_Bits_16___Out_Bits_1___inst0__west_O_layer1_0[0:0];

  assign CB_10_1_inst1__I_6[0:0] = SB_Out_Bits_16___Out_Bits_1___inst0__west_O_layer1_1[0:0];

  assign CB_10_1_inst1__I_7[0:0] = SB_Out_Bits_16___Out_Bits_1___inst0__west_O_layer1_2[0:0];

  assign CB_10_1_inst1__I_8[0:0] = SB_Out_Bits_16___Out_Bits_1___inst0__west_O_layer1_3[0:0];

  assign CB_10_1_inst1__I_9[0:0] = SB_Out_Bits_16___Out_Bits_1___inst0__west_O_layer1_4[0:0];

  assign PECore_inst0__bit1[0:0] = CB_10_1_inst1__O[0:0];

  assign CB_10_1_inst1__clk = clk;

  assign CB_10_1_inst1__config_config_addr[0] = config_config_addr[24];

  assign CB_10_1_inst1__config_config_addr[1] = config_config_addr[25];

  assign CB_10_1_inst1__config_config_addr[2] = config_config_addr[26];

  assign CB_10_1_inst1__config_config_addr[3] = config_config_addr[27];

  assign CB_10_1_inst1__config_config_addr[4] = config_config_addr[28];

  assign CB_10_1_inst1__config_config_addr[5] = config_config_addr[29];

  assign CB_10_1_inst1__config_config_addr[6] = config_config_addr[30];

  assign CB_10_1_inst1__config_config_addr[7] = config_config_addr[31];

  assign CB_10_1_inst1__config_config_data[31:0] = config_config_data[31:0];

  assign CB_10_1_inst1__config_read[0:0] = config_read[0:0];

  assign CB_10_1_inst1__config_write[0] = and_inst7__out;

  assign MuxWithDefaultWrapper_7_32_8_0_inst0__I_5[31:0] = CB_10_1_inst1__read_config_data[31:0];

  assign CB_10_1_inst1__reset = reset;

  assign CB_10_1_inst2__I_0[0:0] = north_I_layer1_0[0:0];

  assign CB_10_1_inst2__I_1[0:0] = north_I_layer1_1[0:0];

  assign CB_10_1_inst2__I_2[0:0] = north_I_layer1_2[0:0];

  assign CB_10_1_inst2__I_3[0:0] = north_I_layer1_3[0:0];

  assign CB_10_1_inst2__I_4[0:0] = north_I_layer1_4[0:0];

  assign CB_10_1_inst2__I_5[0:0] = SB_Out_Bits_16___Out_Bits_1___inst0__north_O_layer1_0[0:0];

  assign CB_10_1_inst2__I_6[0:0] = SB_Out_Bits_16___Out_Bits_1___inst0__north_O_layer1_1[0:0];

  assign CB_10_1_inst2__I_7[0:0] = SB_Out_Bits_16___Out_Bits_1___inst0__north_O_layer1_2[0:0];

  assign CB_10_1_inst2__I_8[0:0] = SB_Out_Bits_16___Out_Bits_1___inst0__north_O_layer1_3[0:0];

  assign CB_10_1_inst2__I_9[0:0] = SB_Out_Bits_16___Out_Bits_1___inst0__north_O_layer1_4[0:0];

  assign PECore_inst0__bit2[0:0] = CB_10_1_inst2__O[0:0];

  assign CB_10_1_inst2__clk = clk;

  assign CB_10_1_inst2__config_config_addr[0] = config_config_addr[24];

  assign CB_10_1_inst2__config_config_addr[1] = config_config_addr[25];

  assign CB_10_1_inst2__config_config_addr[2] = config_config_addr[26];

  assign CB_10_1_inst2__config_config_addr[3] = config_config_addr[27];

  assign CB_10_1_inst2__config_config_addr[4] = config_config_addr[28];

  assign CB_10_1_inst2__config_config_addr[5] = config_config_addr[29];

  assign CB_10_1_inst2__config_config_addr[6] = config_config_addr[30];

  assign CB_10_1_inst2__config_config_addr[7] = config_config_addr[31];

  assign CB_10_1_inst2__config_config_data[31:0] = config_config_data[31:0];

  assign CB_10_1_inst2__config_read[0:0] = config_read[0:0];

  assign CB_10_1_inst2__config_write[0] = and_inst8__out;

  assign MuxWithDefaultWrapper_7_32_8_0_inst0__I_6[31:0] = CB_10_1_inst2__read_config_data[31:0];

  assign CB_10_1_inst2__reset = reset;

  assign Decode08_inst0__I[0] = config_config_addr[16];

  assign Decode08_inst0__I[1] = config_config_addr[17];

  assign Decode08_inst0__I[2] = config_config_addr[18];

  assign Decode08_inst0__I[3] = config_config_addr[19];

  assign Decode08_inst0__I[4] = config_config_addr[20];

  assign Decode08_inst0__I[5] = config_config_addr[21];

  assign Decode08_inst0__I[6] = config_config_addr[22];

  assign Decode08_inst0__I[7] = config_config_addr[23];

  assign and_inst2__in0 = Decode08_inst0__O;

  assign Decode18_inst0__I[0] = config_config_addr[16];

  assign Decode18_inst0__I[1] = config_config_addr[17];

  assign Decode18_inst0__I[2] = config_config_addr[18];

  assign Decode18_inst0__I[3] = config_config_addr[19];

  assign Decode18_inst0__I[4] = config_config_addr[20];

  assign Decode18_inst0__I[5] = config_config_addr[21];

  assign Decode18_inst0__I[6] = config_config_addr[22];

  assign Decode18_inst0__I[7] = config_config_addr[23];

  assign and_inst3__in0 = Decode18_inst0__O;

  assign Decode28_inst0__I[0] = config_config_addr[16];

  assign Decode28_inst0__I[1] = config_config_addr[17];

  assign Decode28_inst0__I[2] = config_config_addr[18];

  assign Decode28_inst0__I[3] = config_config_addr[19];

  assign Decode28_inst0__I[4] = config_config_addr[20];

  assign Decode28_inst0__I[5] = config_config_addr[21];

  assign Decode28_inst0__I[6] = config_config_addr[22];

  assign Decode28_inst0__I[7] = config_config_addr[23];

  assign and_inst4__in0 = Decode28_inst0__O;

  assign Decode38_inst0__I[0] = config_config_addr[16];

  assign Decode38_inst0__I[1] = config_config_addr[17];

  assign Decode38_inst0__I[2] = config_config_addr[18];

  assign Decode38_inst0__I[3] = config_config_addr[19];

  assign Decode38_inst0__I[4] = config_config_addr[20];

  assign Decode38_inst0__I[5] = config_config_addr[21];

  assign Decode38_inst0__I[6] = config_config_addr[22];

  assign Decode38_inst0__I[7] = config_config_addr[23];

  assign and_inst5__in0 = Decode38_inst0__O;

  assign Decode48_inst0__I[0] = config_config_addr[16];

  assign Decode48_inst0__I[1] = config_config_addr[17];

  assign Decode48_inst0__I[2] = config_config_addr[18];

  assign Decode48_inst0__I[3] = config_config_addr[19];

  assign Decode48_inst0__I[4] = config_config_addr[20];

  assign Decode48_inst0__I[5] = config_config_addr[21];

  assign Decode48_inst0__I[6] = config_config_addr[22];

  assign Decode48_inst0__I[7] = config_config_addr[23];

  assign and_inst6__in0 = Decode48_inst0__O;

  assign Decode58_inst0__I[0] = config_config_addr[16];

  assign Decode58_inst0__I[1] = config_config_addr[17];

  assign Decode58_inst0__I[2] = config_config_addr[18];

  assign Decode58_inst0__I[3] = config_config_addr[19];

  assign Decode58_inst0__I[4] = config_config_addr[20];

  assign Decode58_inst0__I[5] = config_config_addr[21];

  assign Decode58_inst0__I[6] = config_config_addr[22];

  assign Decode58_inst0__I[7] = config_config_addr[23];

  assign and_inst7__in0 = Decode58_inst0__O;

  assign Decode68_inst0__I[0] = config_config_addr[16];

  assign Decode68_inst0__I[1] = config_config_addr[17];

  assign Decode68_inst0__I[2] = config_config_addr[18];

  assign Decode68_inst0__I[3] = config_config_addr[19];

  assign Decode68_inst0__I[4] = config_config_addr[20];

  assign Decode68_inst0__I[5] = config_config_addr[21];

  assign Decode68_inst0__I[6] = config_config_addr[22];

  assign Decode68_inst0__I[7] = config_config_addr[23];

  assign and_inst8__in0 = Decode68_inst0__O;

  assign MuxWithDefaultWrapper_7_32_8_0_inst0__EN[0] = and_inst0__out;

  assign MuxWithDefaultWrapper_7_32_8_0_inst0__I_0[31:0] = PECore_inst0__read_config_data[31:0];

  assign MuxWithDefaultWrapper_7_32_8_0_inst0__I_1[31:0] = SB_Out_Bits_16___Out_Bits_1___inst0__read_config_data[31:0];

  assign read_config_data[31:0] = MuxWithDefaultWrapper_7_32_8_0_inst0__O[31:0];

  assign MuxWithDefaultWrapper_7_32_8_0_inst0__S[0] = config_config_addr[16];

  assign MuxWithDefaultWrapper_7_32_8_0_inst0__S[1] = config_config_addr[17];

  assign MuxWithDefaultWrapper_7_32_8_0_inst0__S[2] = config_config_addr[18];

  assign MuxWithDefaultWrapper_7_32_8_0_inst0__S[3] = config_config_addr[19];

  assign MuxWithDefaultWrapper_7_32_8_0_inst0__S[4] = config_config_addr[20];

  assign MuxWithDefaultWrapper_7_32_8_0_inst0__S[5] = config_config_addr[21];

  assign MuxWithDefaultWrapper_7_32_8_0_inst0__S[6] = config_config_addr[22];

  assign MuxWithDefaultWrapper_7_32_8_0_inst0__S[7] = config_config_addr[23];

  assign PECore_inst0__clk = clk;

  assign PECore_inst0__config_config_addr[0] = config_config_addr[24];

  assign PECore_inst0__config_config_addr[1] = config_config_addr[25];

  assign PECore_inst0__config_config_addr[2] = config_config_addr[26];

  assign PECore_inst0__config_config_addr[3] = config_config_addr[27];

  assign PECore_inst0__config_config_addr[4] = config_config_addr[28];

  assign PECore_inst0__config_config_addr[5] = config_config_addr[29];

  assign PECore_inst0__config_config_addr[6] = config_config_addr[30];

  assign PECore_inst0__config_config_addr[7] = config_config_addr[31];

  assign PECore_inst0__config_config_data[31:0] = config_config_data[31:0];

  assign PECore_inst0__config_read[0:0] = config_read[0:0];

  assign PECore_inst0__config_write[0] = and_inst2__out;

  assign SB_Out_Bits_16___Out_Bits_1___inst0__res[15:0] = PECore_inst0__res[15:0];

  assign SB_Out_Bits_16___Out_Bits_1___inst0__res_p[0:0] = PECore_inst0__res_p[0:0];

  assign PECore_inst0__reset = reset;

  assign PECore_inst0__stall[3:0] = stall[3:0];

  assign SB_Out_Bits_16___Out_Bits_1___inst0__clk = clk;

  assign SB_Out_Bits_16___Out_Bits_1___inst0__config_config_addr[0] = config_config_addr[24];

  assign SB_Out_Bits_16___Out_Bits_1___inst0__config_config_addr[1] = config_config_addr[25];

  assign SB_Out_Bits_16___Out_Bits_1___inst0__config_config_addr[2] = config_config_addr[26];

  assign SB_Out_Bits_16___Out_Bits_1___inst0__config_config_addr[3] = config_config_addr[27];

  assign SB_Out_Bits_16___Out_Bits_1___inst0__config_config_addr[4] = config_config_addr[28];

  assign SB_Out_Bits_16___Out_Bits_1___inst0__config_config_addr[5] = config_config_addr[29];

  assign SB_Out_Bits_16___Out_Bits_1___inst0__config_config_addr[6] = config_config_addr[30];

  assign SB_Out_Bits_16___Out_Bits_1___inst0__config_config_addr[7] = config_config_addr[31];

  assign SB_Out_Bits_16___Out_Bits_1___inst0__config_config_data[31:0] = config_config_data[31:0];

  assign SB_Out_Bits_16___Out_Bits_1___inst0__config_read[0:0] = config_read[0:0];

  assign SB_Out_Bits_16___Out_Bits_1___inst0__config_write[0] = and_inst3__out;

  assign SB_Out_Bits_16___Out_Bits_1___inst0__east_I_layer16_0[15:0] = east_I_layer16_0[15:0];

  assign SB_Out_Bits_16___Out_Bits_1___inst0__east_I_layer16_1[15:0] = east_I_layer16_1[15:0];

  assign SB_Out_Bits_16___Out_Bits_1___inst0__east_I_layer16_2[15:0] = east_I_layer16_2[15:0];

  assign SB_Out_Bits_16___Out_Bits_1___inst0__east_I_layer16_3[15:0] = east_I_layer16_3[15:0];

  assign SB_Out_Bits_16___Out_Bits_1___inst0__east_I_layer16_4[15:0] = east_I_layer16_4[15:0];

  assign SB_Out_Bits_16___Out_Bits_1___inst0__east_I_layer1_0[0:0] = east_I_layer1_0[0:0];

  assign SB_Out_Bits_16___Out_Bits_1___inst0__east_I_layer1_1[0:0] = east_I_layer1_1[0:0];

  assign SB_Out_Bits_16___Out_Bits_1___inst0__east_I_layer1_2[0:0] = east_I_layer1_2[0:0];

  assign SB_Out_Bits_16___Out_Bits_1___inst0__east_I_layer1_3[0:0] = east_I_layer1_3[0:0];

  assign SB_Out_Bits_16___Out_Bits_1___inst0__east_I_layer1_4[0:0] = east_I_layer1_4[0:0];

  assign east_O_layer16_0[15:0] = SB_Out_Bits_16___Out_Bits_1___inst0__east_O_layer16_0[15:0];

  assign east_O_layer16_1[15:0] = SB_Out_Bits_16___Out_Bits_1___inst0__east_O_layer16_1[15:0];

  assign east_O_layer16_2[15:0] = SB_Out_Bits_16___Out_Bits_1___inst0__east_O_layer16_2[15:0];

  assign east_O_layer16_3[15:0] = SB_Out_Bits_16___Out_Bits_1___inst0__east_O_layer16_3[15:0];

  assign east_O_layer16_4[15:0] = SB_Out_Bits_16___Out_Bits_1___inst0__east_O_layer16_4[15:0];

  assign east_O_layer1_0[0:0] = SB_Out_Bits_16___Out_Bits_1___inst0__east_O_layer1_0[0:0];

  assign east_O_layer1_1[0:0] = SB_Out_Bits_16___Out_Bits_1___inst0__east_O_layer1_1[0:0];

  assign east_O_layer1_2[0:0] = SB_Out_Bits_16___Out_Bits_1___inst0__east_O_layer1_2[0:0];

  assign east_O_layer1_3[0:0] = SB_Out_Bits_16___Out_Bits_1___inst0__east_O_layer1_3[0:0];

  assign east_O_layer1_4[0:0] = SB_Out_Bits_16___Out_Bits_1___inst0__east_O_layer1_4[0:0];

  assign SB_Out_Bits_16___Out_Bits_1___inst0__north_I_layer16_0[15:0] = north_I_layer16_0[15:0];

  assign SB_Out_Bits_16___Out_Bits_1___inst0__north_I_layer16_1[15:0] = north_I_layer16_1[15:0];

  assign SB_Out_Bits_16___Out_Bits_1___inst0__north_I_layer16_2[15:0] = north_I_layer16_2[15:0];

  assign SB_Out_Bits_16___Out_Bits_1___inst0__north_I_layer16_3[15:0] = north_I_layer16_3[15:0];

  assign SB_Out_Bits_16___Out_Bits_1___inst0__north_I_layer16_4[15:0] = north_I_layer16_4[15:0];

  assign SB_Out_Bits_16___Out_Bits_1___inst0__north_I_layer1_0[0:0] = north_I_layer1_0[0:0];

  assign SB_Out_Bits_16___Out_Bits_1___inst0__north_I_layer1_1[0:0] = north_I_layer1_1[0:0];

  assign SB_Out_Bits_16___Out_Bits_1___inst0__north_I_layer1_2[0:0] = north_I_layer1_2[0:0];

  assign SB_Out_Bits_16___Out_Bits_1___inst0__north_I_layer1_3[0:0] = north_I_layer1_3[0:0];

  assign SB_Out_Bits_16___Out_Bits_1___inst0__north_I_layer1_4[0:0] = north_I_layer1_4[0:0];

  assign north_O_layer16_0[15:0] = SB_Out_Bits_16___Out_Bits_1___inst0__north_O_layer16_0[15:0];

  assign north_O_layer16_1[15:0] = SB_Out_Bits_16___Out_Bits_1___inst0__north_O_layer16_1[15:0];

  assign north_O_layer16_2[15:0] = SB_Out_Bits_16___Out_Bits_1___inst0__north_O_layer16_2[15:0];

  assign north_O_layer16_3[15:0] = SB_Out_Bits_16___Out_Bits_1___inst0__north_O_layer16_3[15:0];

  assign north_O_layer16_4[15:0] = SB_Out_Bits_16___Out_Bits_1___inst0__north_O_layer16_4[15:0];

  assign north_O_layer1_0[0:0] = SB_Out_Bits_16___Out_Bits_1___inst0__north_O_layer1_0[0:0];

  assign north_O_layer1_1[0:0] = SB_Out_Bits_16___Out_Bits_1___inst0__north_O_layer1_1[0:0];

  assign north_O_layer1_2[0:0] = SB_Out_Bits_16___Out_Bits_1___inst0__north_O_layer1_2[0:0];

  assign north_O_layer1_3[0:0] = SB_Out_Bits_16___Out_Bits_1___inst0__north_O_layer1_3[0:0];

  assign north_O_layer1_4[0:0] = SB_Out_Bits_16___Out_Bits_1___inst0__north_O_layer1_4[0:0];

  assign SB_Out_Bits_16___Out_Bits_1___inst0__reset = reset;

  assign SB_Out_Bits_16___Out_Bits_1___inst0__south_I_layer16_0[15:0] = south_I_layer16_0[15:0];

  assign SB_Out_Bits_16___Out_Bits_1___inst0__south_I_layer16_1[15:0] = south_I_layer16_1[15:0];

  assign SB_Out_Bits_16___Out_Bits_1___inst0__south_I_layer16_2[15:0] = south_I_layer16_2[15:0];

  assign SB_Out_Bits_16___Out_Bits_1___inst0__south_I_layer16_3[15:0] = south_I_layer16_3[15:0];

  assign SB_Out_Bits_16___Out_Bits_1___inst0__south_I_layer16_4[15:0] = south_I_layer16_4[15:0];

  assign SB_Out_Bits_16___Out_Bits_1___inst0__south_I_layer1_0[0:0] = south_I_layer1_0[0:0];

  assign SB_Out_Bits_16___Out_Bits_1___inst0__south_I_layer1_1[0:0] = south_I_layer1_1[0:0];

  assign SB_Out_Bits_16___Out_Bits_1___inst0__south_I_layer1_2[0:0] = south_I_layer1_2[0:0];

  assign SB_Out_Bits_16___Out_Bits_1___inst0__south_I_layer1_3[0:0] = south_I_layer1_3[0:0];

  assign SB_Out_Bits_16___Out_Bits_1___inst0__south_I_layer1_4[0:0] = south_I_layer1_4[0:0];

  assign south_O_layer16_0[15:0] = SB_Out_Bits_16___Out_Bits_1___inst0__south_O_layer16_0[15:0];

  assign south_O_layer16_1[15:0] = SB_Out_Bits_16___Out_Bits_1___inst0__south_O_layer16_1[15:0];

  assign south_O_layer16_2[15:0] = SB_Out_Bits_16___Out_Bits_1___inst0__south_O_layer16_2[15:0];

  assign south_O_layer16_3[15:0] = SB_Out_Bits_16___Out_Bits_1___inst0__south_O_layer16_3[15:0];

  assign south_O_layer16_4[15:0] = SB_Out_Bits_16___Out_Bits_1___inst0__south_O_layer16_4[15:0];

  assign south_O_layer1_0[0:0] = SB_Out_Bits_16___Out_Bits_1___inst0__south_O_layer1_0[0:0];

  assign south_O_layer1_1[0:0] = SB_Out_Bits_16___Out_Bits_1___inst0__south_O_layer1_1[0:0];

  assign south_O_layer1_2[0:0] = SB_Out_Bits_16___Out_Bits_1___inst0__south_O_layer1_2[0:0];

  assign south_O_layer1_3[0:0] = SB_Out_Bits_16___Out_Bits_1___inst0__south_O_layer1_3[0:0];

  assign south_O_layer1_4[0:0] = SB_Out_Bits_16___Out_Bits_1___inst0__south_O_layer1_4[0:0];

  assign SB_Out_Bits_16___Out_Bits_1___inst0__west_I_layer16_0[15:0] = west_I_layer16_0[15:0];

  assign SB_Out_Bits_16___Out_Bits_1___inst0__west_I_layer16_1[15:0] = west_I_layer16_1[15:0];

  assign SB_Out_Bits_16___Out_Bits_1___inst0__west_I_layer16_2[15:0] = west_I_layer16_2[15:0];

  assign SB_Out_Bits_16___Out_Bits_1___inst0__west_I_layer16_3[15:0] = west_I_layer16_3[15:0];

  assign SB_Out_Bits_16___Out_Bits_1___inst0__west_I_layer16_4[15:0] = west_I_layer16_4[15:0];

  assign SB_Out_Bits_16___Out_Bits_1___inst0__west_I_layer1_0[0:0] = west_I_layer1_0[0:0];

  assign SB_Out_Bits_16___Out_Bits_1___inst0__west_I_layer1_1[0:0] = west_I_layer1_1[0:0];

  assign SB_Out_Bits_16___Out_Bits_1___inst0__west_I_layer1_2[0:0] = west_I_layer1_2[0:0];

  assign SB_Out_Bits_16___Out_Bits_1___inst0__west_I_layer1_3[0:0] = west_I_layer1_3[0:0];

  assign SB_Out_Bits_16___Out_Bits_1___inst0__west_I_layer1_4[0:0] = west_I_layer1_4[0:0];

  assign west_O_layer16_0[15:0] = SB_Out_Bits_16___Out_Bits_1___inst0__west_O_layer16_0[15:0];

  assign west_O_layer16_1[15:0] = SB_Out_Bits_16___Out_Bits_1___inst0__west_O_layer16_1[15:0];

  assign west_O_layer16_2[15:0] = SB_Out_Bits_16___Out_Bits_1___inst0__west_O_layer16_2[15:0];

  assign west_O_layer16_3[15:0] = SB_Out_Bits_16___Out_Bits_1___inst0__west_O_layer16_3[15:0];

  assign west_O_layer16_4[15:0] = SB_Out_Bits_16___Out_Bits_1___inst0__west_O_layer16_4[15:0];

  assign west_O_layer1_0[0:0] = SB_Out_Bits_16___Out_Bits_1___inst0__west_O_layer1_0[0:0];

  assign west_O_layer1_1[0:0] = SB_Out_Bits_16___Out_Bits_1___inst0__west_O_layer1_1[0:0];

  assign west_O_layer1_2[0:0] = SB_Out_Bits_16___Out_Bits_1___inst0__west_O_layer1_2[0:0];

  assign west_O_layer1_3[0:0] = SB_Out_Bits_16___Out_Bits_1___inst0__west_O_layer1_3[0:0];

  assign west_O_layer1_4[0:0] = SB_Out_Bits_16___Out_Bits_1___inst0__west_O_layer1_4[0:0];

  assign and_inst0__in0 = coreir_eq_16_inst0__out;

  assign and_inst0__in1 = config_read[0];

  assign and_inst1__in0 = coreir_eq_16_inst0__out;

  assign and_inst1__in1 = config_write[0];

  assign and_inst2__in1 = and_inst1__out;

  assign and_inst3__in1 = and_inst1__out;

  assign and_inst4__in1 = and_inst1__out;

  assign and_inst5__in1 = and_inst1__out;

  assign and_inst6__in1 = and_inst1__out;

  assign and_inst7__in1 = and_inst1__out;

  assign and_inst8__in1 = and_inst1__out;

  assign coreir_eq_16_inst0__in0[15:0] = tile_id[15:0];

  assign coreir_eq_16_inst0__in1[0] = config_config_addr[0];

  assign coreir_eq_16_inst0__in1[10] = config_config_addr[10];

  assign coreir_eq_16_inst0__in1[11] = config_config_addr[11];

  assign coreir_eq_16_inst0__in1[12] = config_config_addr[12];

  assign coreir_eq_16_inst0__in1[13] = config_config_addr[13];

  assign coreir_eq_16_inst0__in1[14] = config_config_addr[14];

  assign coreir_eq_16_inst0__in1[15] = config_config_addr[15];

  assign coreir_eq_16_inst0__in1[1] = config_config_addr[1];

  assign coreir_eq_16_inst0__in1[2] = config_config_addr[2];

  assign coreir_eq_16_inst0__in1[3] = config_config_addr[3];

  assign coreir_eq_16_inst0__in1[4] = config_config_addr[4];

  assign coreir_eq_16_inst0__in1[5] = config_config_addr[5];

  assign coreir_eq_16_inst0__in1[6] = config_config_addr[6];

  assign coreir_eq_16_inst0__in1[7] = config_config_addr[7];

  assign coreir_eq_16_inst0__in1[8] = config_config_addr[8];

  assign coreir_eq_16_inst0__in1[9] = config_config_addr[9];


endmodule  // Tile_PECore

